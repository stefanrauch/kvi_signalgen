flash_loader_inst : flash_loader PORT MAP (
		noe_in	 => noe_in_sig
	);
