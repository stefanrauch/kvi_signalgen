-- megafunction wizard: %ALTASMI_PARALLEL%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: ALTASMI_PARALLEL 

-- ============================================================
-- File Name: flash_access.vhd
-- Megafunction Name(s):
-- 			ALTASMI_PARALLEL
--
-- Simulation Library Files(s):
-- 			
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 11.1 Build 173 11/01/2011 SJ Full Version
-- ************************************************************


--Copyright (C) 1991-2011 Altera Corporation
--Your use of Altera Corporation's design tools, logic functions 
--and other software and tools, and its AMPP partner logic 
--functions, and any output files from any of the foregoing 
--(including device programming or simulation files), and any 
--associated documentation or information are expressly subject 
--to the terms and conditions of the Altera Program License 
--Subscription Agreement, Altera MegaCore Function License 
--Agreement, or other applicable license agreement, including, 
--without limitation, that your use is for the sole purpose of 
--programming logic devices manufactured by Altera and sold by 
--Altera or its authorized distributors.  Please refer to the 
--applicable agreement for further details.


--altasmi_parallel CBX_AUTO_BLACKBOX="ALL" DATA_WIDTH="STANDARD" DEVICE_FAMILY="Arria II GX" EPCS_TYPE="EPCS128" PAGE_SIZE=256 PORT_BULK_ERASE="PORT_UNUSED" PORT_FAST_READ="PORT_UNUSED" PORT_ILLEGAL_ERASE="PORT_USED" PORT_ILLEGAL_WRITE="PORT_USED" PORT_RDID_OUT="PORT_USED" PORT_READ_ADDRESS="PORT_UNUSED" PORT_READ_RDID="PORT_USED" PORT_READ_SID="PORT_UNUSED" PORT_READ_STATUS="PORT_USED" PORT_SECTOR_ERASE="PORT_USED" PORT_SECTOR_PROTECT="PORT_UNUSED" PORT_SHIFT_BYTES="PORT_USED" PORT_WREN="PORT_USED" PORT_WRITE="PORT_USED" USE_EAB="ON" addr busy clkin data_valid datain dataout illegal_erase illegal_write rden rdid_out read read_rdid read_status sector_erase shift_bytes status_out wren write INTENDED_DEVICE_FAMILY="Arria II GX" ALTERA_INTERNAL_OPTIONS=SUPPRESS_DA_RULE_INTERNAL=C106
--VERSION_BEGIN 11.1 cbx_a_gray2bin 2011:10:31:21:13:12:SJ cbx_a_graycounter 2011:10:31:21:13:12:SJ cbx_altasmi_parallel 2011:10:31:21:13:12:SJ cbx_altdpram 2011:10:31:21:13:12:SJ cbx_altsyncram 2011:10:31:21:13:13:SJ cbx_cyclone 2011:10:31:21:13:13:SJ cbx_cycloneii 2011:10:31:21:13:13:SJ cbx_fifo_common 2011:10:31:21:13:12:SJ cbx_lpm_add_sub 2011:10:31:21:13:13:SJ cbx_lpm_compare 2011:10:31:21:13:13:SJ cbx_lpm_counter 2011:10:31:21:13:13:SJ cbx_lpm_decode 2011:10:31:21:13:13:SJ cbx_lpm_mux 2011:10:31:21:13:13:SJ cbx_mgl 2011:10:31:21:15:34:SJ cbx_scfifo 2011:10:31:21:13:14:SJ cbx_stratix 2011:10:31:21:13:14:SJ cbx_stratixii 2011:10:31:21:13:14:SJ cbx_stratixiii 2011:10:31:21:13:14:SJ cbx_stratixv 2011:10:31:21:13:14:SJ cbx_util_mgl 2011:10:31:21:13:14:SJ  VERSION_END

 LIBRARY altera_mf;
 USE altera_mf.all;

 LIBRARY arriaii;
 USE arriaii.all;

 LIBRARY lpm;
 USE lpm.all;

--synthesis_resources = a_graycounter 4 arriaii_asmiblock 1 lpm_compare 2 lpm_counter 2 lut 29 mux21 1 reg 126 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  flash_access_altasmi_parallel_era2 IS 
	 PORT 
	 ( 
		 addr	:	IN  STD_LOGIC_VECTOR (23 DOWNTO 0);
		 busy	:	OUT  STD_LOGIC;
		 clkin	:	IN  STD_LOGIC;
		 data_valid	:	OUT  STD_LOGIC;
		 datain	:	IN  STD_LOGIC_VECTOR (7 DOWNTO 0) := (OTHERS => '0');
		 dataout	:	OUT  STD_LOGIC_VECTOR (7 DOWNTO 0);
		 illegal_erase	:	OUT  STD_LOGIC;
		 illegal_write	:	OUT  STD_LOGIC;
		 rden	:	IN  STD_LOGIC;
		 rdid_out	:	OUT  STD_LOGIC_VECTOR (7 DOWNTO 0);
		 read	:	IN  STD_LOGIC := '0';
		 read_rdid	:	IN  STD_LOGIC := '0';
		 read_status	:	IN  STD_LOGIC := '0';
		 sector_erase	:	IN  STD_LOGIC := '0';
		 shift_bytes	:	IN  STD_LOGIC := '0';
		 status_out	:	OUT  STD_LOGIC_VECTOR (7 DOWNTO 0);
		 wren	:	IN  STD_LOGIC := '1';
		 write	:	IN  STD_LOGIC := '0'
	 ); 
 END flash_access_altasmi_parallel_era2;

 ARCHITECTURE RTL OF flash_access_altasmi_parallel_era2 IS

	 ATTRIBUTE synthesis_clearbox : natural;
	 ATTRIBUTE synthesis_clearbox OF RTL : ARCHITECTURE IS 2;
	 ATTRIBUTE ALTERA_ATTRIBUTE : string;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF RTL : ARCHITECTURE IS "SUPPRESS_DA_RULE_INTERNAL=C106";

	 SIGNAL  wire_addbyte_cntr_w_lg_w_q_range123w124w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_addbyte_cntr_w_lg_w_q_range121w122w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_addbyte_cntr_clk_en	:	STD_LOGIC;
	 SIGNAL  wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range82w85w118w119w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_addbyte_cntr_clock	:	STD_LOGIC;
	 SIGNAL  wire_addbyte_cntr_q	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_addbyte_cntr_w_q_range121w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_addbyte_cntr_w_q_range123w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_gen_cntr_w_lg_w_q_range92w93w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_gen_cntr_w_lg_w_q_range90w91w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_gen_cntr_clk_en	:	STD_LOGIC;
	 SIGNAL  wire_w_lg_in_operation36w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_gen_cntr_q	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_gen_cntr_w_q_range90w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_gen_cntr_w_q_range92w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w220w221w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w220w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w225w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_lg_w_lg_w_lg_w_q_range82w85w217w218w219w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_lg_w_lg_w_lg_w_q_range82w85w222w223w224w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_lg_w_lg_w_lg_w_q_range82w83w84w229w230w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range82w87w293w294w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range82w85w234w235w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range82w85w240w241w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range82w85w217w218w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range82w85w222w223w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range82w83w84w229w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_lg_w_q_range82w87w293w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_lg_w_q_range82w85w234w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_lg_w_q_range82w85w240w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_lg_w_q_range82w85w217w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_lg_w_q_range82w85w222w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_lg_w_q_range82w85w118w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_lg_w_lg_w_lg_w_q_range81w86w100w101w102w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_lg_w_q_range81w86w100w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_lg_w_q_range82w83w84w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_q_range82w87w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_q_range82w85w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range81w86w100w101w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_q_range81w86w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_q_range82w83w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_clk_en	:	STD_LOGIC;
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_w_lg_w74w75w76w77w78w79w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_q	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_q_range81w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_q_range82w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_wrstage_cntr_w_lg_w_q_range462w463w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_wrstage_cntr_w_lg_w_q_range460w461w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_wrstage_cntr_clk_en	:	STD_LOGIC;
	 SIGNAL  wire_w459w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_wrstage_cntr_clock	:	STD_LOGIC;
	 SIGNAL  wire_wrstage_cntr_q	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_wrstage_cntr_w_q_range460w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_wrstage_cntr_w_q_range462w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 add_msb_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_add_msb_reg_ena	:	STD_LOGIC;
	 SIGNAL	 wire_addr_reg_d	:	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL	 addr_reg	:	STD_LOGIC_VECTOR(23 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_addr_reg_ena	:	STD_LOGIC_VECTOR(23 DOWNTO 0);
	 SIGNAL  wire_addr_reg_w_lg_w_lg_w_lg_w506w507w508w509w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_addr_reg_w_lg_w_lg_w506w507w508w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_addr_reg_w_lg_w498w499w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_addr_reg_w_lg_w502w503w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_addr_reg_w_lg_w506w507w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_addr_reg_w498w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_addr_reg_w502w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_addr_reg_w506w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_addr_reg_w_lg_w_lg_w_lg_w_lg_w_q_range297w485w486w487w488w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_addr_reg_w_lg_w_lg_w_lg_w_lg_w_q_range297w485w490w496w497w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_addr_reg_w_lg_w_lg_w_lg_w_lg_w_q_range297w485w490w496w501w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_addr_reg_w_lg_w_lg_w_lg_w_q_range297w485w486w487w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_addr_reg_w_lg_w_lg_w_lg_w_q_range297w485w490w491w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_addr_reg_w_lg_w_lg_w_lg_w_q_range297w485w490w496w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_addr_reg_w_lg_w_lg_w_q_range297w480w481w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_addr_reg_w_lg_w_lg_w_q_range297w485w486w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_addr_reg_w_lg_w_lg_w_q_range297w485w490w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_addr_reg_w_lg_w_q_range297w480w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_addr_reg_w_lg_w_q_range297w485w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_addr_reg_w_q_range505w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_addr_reg_w_q_range500w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_addr_reg_w_q_range495w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_addr_reg_w_q_range489w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_addr_reg_w_q_range272w	:	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  wire_addr_reg_w_q_range484w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_addr_reg_w_q_range297w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 wire_asmi_opcode_reg_d	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL	 asmi_opcode_reg	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_asmi_opcode_reg_ena	:	STD_LOGIC_VECTOR(7 DOWNTO 0);
	 SIGNAL  wire_asmi_opcode_reg_w_q_range129w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL	 buf_empty_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 busy_det_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 clr_addmsb_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 clr_endrbyte_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_clr_endrbyte_reg_w_lg_q359w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 clr_rdid_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 clr_rdid_reg2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 clr_read_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 clr_read_reg2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 clr_rstat_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 clr_rstat_reg2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 clr_write_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 clr_write_reg2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 cnt_bfend_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 do_wrmemadd_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 dvalid_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_dvalid_reg_ena	:	STD_LOGIC;
	 SIGNAL	 dvalid_reg2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 end1_cyc_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 end1_cyc_reg2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 end_op_hdlyreg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 end_op_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 end_pgwrop_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_end_pgwrop_reg_ena	:	STD_LOGIC;
	 SIGNAL	 end_rbyte_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_end_rbyte_reg_ena	:	STD_LOGIC;
	 SIGNAL	 end_read_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 ill_erase_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 ill_write_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 max_cnt_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 maxcnt_shift_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 maxcnt_shift_reg2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 ncs_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_ncs_reg_ena	:	STD_LOGIC;
	 SIGNAL  wire_ncs_reg_w_lg_q262w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 wire_pgwrbuf_dataout_d	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL	 pgwrbuf_dataout	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_pgwrbuf_dataout_ena	:	STD_LOGIC_VECTOR(7 DOWNTO 0);
	 SIGNAL  wire_pgwrbuf_dataout_w_q_range407w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL	 rdid_out_reg	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 read_bufdly_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_read_data_reg_d	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL	 read_data_reg	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_read_data_reg_ena	:	STD_LOGIC_VECTOR(7 DOWNTO 0);
	 SIGNAL	 wire_read_dout_reg_d	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL	 read_dout_reg	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_read_dout_reg_ena	:	STD_LOGIC_VECTOR(7 DOWNTO 0);
	 SIGNAL	 read_rdid_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 read_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_read_reg_ena	:	STD_LOGIC;
	 SIGNAL	 read_status_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sec_erase_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_sec_erase_reg_ena	:	STD_LOGIC;
	 SIGNAL	 shftpgwr_data_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 shift_op_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 stage2_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 stage3_dly_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 stage3_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 stage4_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 start_wrpoll_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_start_wrpoll_reg_ena	:	STD_LOGIC;
	 SIGNAL	 start_wrpoll_reg2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_statreg_int_d	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL	 statreg_int	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_statreg_int_ena	:	STD_LOGIC_VECTOR(7 DOWNTO 0);
	 SIGNAL	 wire_statreg_out_d	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL	 statreg_out	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_statreg_out_ena	:	STD_LOGIC_VECTOR(7 DOWNTO 0);
	 SIGNAL	 write_prot_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_write_prot_reg_ena	:	STD_LOGIC;
	 SIGNAL	 write_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_write_reg_ena	:	STD_LOGIC;
	 SIGNAL	 write_rstat_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_cmpr4_aeb	:	STD_LOGIC;
	 SIGNAL  wire_cmpr4_dataa	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_cmpr4_datab	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_cmpr5_aeb	:	STD_LOGIC;
	 SIGNAL  wire_cmpr5_dataa	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_cmpr5_datab	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_pgwr_data_cntr_clk_en	:	STD_LOGIC;
	 SIGNAL  wire_w_lg_w_lg_w_lg_shift_bytes_wire403w419w420w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_pgwr_data_cntr_q	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_pgwr_data_cntr_w_q_range424w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_pgwr_data_cntr_w_q_range427w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_pgwr_data_cntr_w_q_range430w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_pgwr_data_cntr_w_q_range433w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_pgwr_data_cntr_w_q_range436w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_pgwr_data_cntr_w_q_range439w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_pgwr_data_cntr_w_q_range442w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_pgwr_data_cntr_w_q_range445w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_pgwr_read_cntr_q	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL	wire_mux211_dataout	:	STD_LOGIC;
	 SIGNAL  wire_scfifo3_data	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_scfifo3_q	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_scfifo3_rdreq	:	STD_LOGIC;
	 SIGNAL  wire_w_lg_read_buf405w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_scfifo3_wrreq	:	STD_LOGIC;
	 SIGNAL  wire_w_lg_w_lg_shift_bytes_wire403w404w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_scfifo3_w_q_range410w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_scfifo3_w_q_range415w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stratixii_asmiblock2_data0out	:	STD_LOGIC;
	 SIGNAL  wire_w383w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w348w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_end_operation379w380w381w382w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_load_opcode135w136w137w184w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_load_opcode135w136w137w138w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_load_opcode140w141w142w186w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_load_opcode140w141w142w143w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_load_opcode159w160w161w196w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_load_opcode159w160w161w162w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_do_read245w246w247w248w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_do_write378w552w553w554w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w555w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_do_read301w345w346w347w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_do_sec_erase289w290w291w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_end_operation379w380w381w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_load_opcode135w136w137w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_load_opcode140w141w142w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_load_opcode159w160w161w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_do_read245w246w247w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_do_read245w246w292w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_do_write378w552w553w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_do_write57w58w548w549w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_do_read301w345w346w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_bp2_wire477w478w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_do_polling389w390w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_do_sec_erase289w290w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_do_write148w149w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_do_write48w226w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_end_operation379w380w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode150w190w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode150w151w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode135w136w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode153w192w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode153w154w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode156w194w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode156w157w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode164w198w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode164w165w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode167w200w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode167w168w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode145w188w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode145w146w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode140w141w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode159w160w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode132w182w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode132w133w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_reach_max_cnt453w454w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_start_poll231w232w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_do_read245w246w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_do_write378w552w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_read_bufdly408w409w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_do_write57w58w457w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_do_write57w58w59w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_do_write57w58w548w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_do_read301w345w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_do_write57w282w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_end_operation391w392w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_rden_wire286w287w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_bp2_wire477w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_bulk_erase227w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_polling389w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_sec_erase289w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_write148w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_write55w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_write48w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_end_operation379w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_load_opcode150w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_load_opcode135w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_load_opcode153w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_load_opcode156w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_load_opcode164w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_load_opcode167w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_load_opcode145w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_load_opcode140w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_load_opcode159w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_load_opcode132w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_not_busy280w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_not_busy275w	:	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  wire_w_lg_reach_max_cnt453w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_bufdly416w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_bufdly411w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_shift_opcode130w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_stage3_wire285w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_stage3_wire312w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_stage3_wire273w	:	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  wire_w_lg_stage4_wire314w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_start_poll231w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_do_write48w243w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_bp0_wire479w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_bp1_wire483w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_bp2_wire494w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_buf_empty524w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_busy_wire1w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_clkin_wire80w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_bulk_erase376w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_fast_read244w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_memadd298w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_polling239w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_read245w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_read_rdid37w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_read_stat38w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_sec_erase377w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_sec_prot375w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_wren39w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_write378w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_end_add_cycle67w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_end_fast_read61w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_end_ophdly35w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_end_pgwr_data47w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_end_read64w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_rden_wire360w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_reach_max_cnt418w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_bufdly408w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_rdid_wire10w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_sid_wire9w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_status_wire23w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_sec_protect_wire8w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_st_busy_wire95w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_prot_true456w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_wire18w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_pagewr_buf_not_empty_range53w54w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w555w556w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_load_opcode167w200w201w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_load_opcode167w168w169w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_do_write57w282w283w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_rden_wire286w287w288w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_not_busy275w276w	:	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_read_bufdly411w412w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_stage4_wire314w315w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_load_opcode167w200w201w202w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_load_opcode167w168w169w170w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_do_write57w282w283w284w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w203w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w171w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w203w204w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w171w172w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w203w204w205w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w171w172w173w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w203w204w205w206w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w171w172w173w174w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_w203w204w205w206w207w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_w171w172w173w174w175w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_w_lg_w203w204w205w206w207w208w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_w_lg_w171w172w173w174w175w176w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w209w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w177w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w177w178w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w117w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_do_read_sid113w114w115w116w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_do_read301w302w303w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_do_read_sid113w114w115w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_do_read301w313w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_do_read301w302w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_do_read_sid113w114w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_do_sec_erase468w469w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_do_write57w58w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_data0out_wire317w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_read301w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_read_sid113w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_read_stat311w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_sec_erase468w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_wren228w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_write57w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_end_operation391w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_load_opcode211w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_rden_wire286w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_bufdly406w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_pagewr_buf_not_empty_range422w425w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_pagewr_buf_not_empty_range426w428w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_pagewr_buf_not_empty_range429w431w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_pagewr_buf_not_empty_range432w434w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_pagewr_buf_not_empty_range435w437w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_pagewr_buf_not_empty_range438w440w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_pagewr_buf_not_empty_range441w443w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_pagewr_buf_not_empty_range444w446w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  be_write_prot :	STD_LOGIC;
	 SIGNAL  berase_opcode :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  bp0_wire :	STD_LOGIC;
	 SIGNAL  bp1_wire :	STD_LOGIC;
	 SIGNAL  bp2_wire :	STD_LOGIC;
	 SIGNAL  bp3_wire :	STD_LOGIC;
	 SIGNAL  buf_empty :	STD_LOGIC;
	 SIGNAL  busy_wire :	STD_LOGIC;
	 SIGNAL  clkin_wire :	STD_LOGIC;
	 SIGNAL  clr_rdid_wire :	STD_LOGIC;
	 SIGNAL  clr_read_wire :	STD_LOGIC;
	 SIGNAL  clr_rstat_wire :	STD_LOGIC;
	 SIGNAL  clr_write_wire :	STD_LOGIC;
	 SIGNAL  cnt_bfend_wire_in :	STD_LOGIC;
	 SIGNAL  data0out_wire :	STD_LOGIC;
	 SIGNAL  data_valid_wire :	STD_LOGIC;
	 SIGNAL  dataout_wire :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  do_bulk_erase :	STD_LOGIC;
	 SIGNAL  do_fast_read :	STD_LOGIC;
	 SIGNAL  do_memadd :	STD_LOGIC;
	 SIGNAL  do_polling :	STD_LOGIC;
	 SIGNAL  do_read :	STD_LOGIC;
	 SIGNAL  do_read_rdid :	STD_LOGIC;
	 SIGNAL  do_read_sid :	STD_LOGIC;
	 SIGNAL  do_read_stat :	STD_LOGIC;
	 SIGNAL  do_sec_erase :	STD_LOGIC;
	 SIGNAL  do_sec_prot :	STD_LOGIC;
	 SIGNAL  do_secprot_wren :	STD_LOGIC;
	 SIGNAL  do_sprot_polling :	STD_LOGIC;
	 SIGNAL  do_sprot_rstat :	STD_LOGIC;
	 SIGNAL  do_wren :	STD_LOGIC;
	 SIGNAL  do_write :	STD_LOGIC;
	 SIGNAL  do_write_polling :	STD_LOGIC;
	 SIGNAL  do_write_rstat :	STD_LOGIC;
	 SIGNAL  do_write_wren :	STD_LOGIC;
	 SIGNAL  dummy_read_buf :	STD_LOGIC;
	 SIGNAL  end1_cyc_gen_cntr_wire :	STD_LOGIC;
	 SIGNAL  end1_cyc_normal_in_wire :	STD_LOGIC;
	 SIGNAL  end1_cyc_reg_in_wire :	STD_LOGIC;
	 SIGNAL  end_add_cycle :	STD_LOGIC;
	 SIGNAL  end_add_cycle_mux_datab_wire :	STD_LOGIC;
	 SIGNAL  end_fast_read :	STD_LOGIC;
	 SIGNAL  end_one_cyc_pos :	STD_LOGIC;
	 SIGNAL  end_one_cycle :	STD_LOGIC;
	 SIGNAL  end_operation :	STD_LOGIC;
	 SIGNAL  end_ophdly :	STD_LOGIC;
	 SIGNAL  end_pgwr_data :	STD_LOGIC;
	 SIGNAL  end_read :	STD_LOGIC;
	 SIGNAL  end_read_byte :	STD_LOGIC;
	 SIGNAL  end_wrstage :	STD_LOGIC;
	 SIGNAL  fast_read_opcode :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  fast_read_wire :	STD_LOGIC;
	 SIGNAL  ill_erase_wire :	STD_LOGIC;
	 SIGNAL  ill_write_wire :	STD_LOGIC;
	 SIGNAL  illegal_erase_b4out_wire :	STD_LOGIC;
	 SIGNAL  illegal_write_b4out_wire :	STD_LOGIC;
	 SIGNAL  in_operation :	STD_LOGIC;
	 SIGNAL  load_opcode :	STD_LOGIC;
	 SIGNAL  memadd_sdoin :	STD_LOGIC;
	 SIGNAL  not_busy :	STD_LOGIC;
	 SIGNAL  oe_wire :	STD_LOGIC;
	 SIGNAL  page_size_wire :	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  pagewr_buf_not_empty :	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  rden_wire :	STD_LOGIC;
	 SIGNAL  rdid_load :	STD_LOGIC;
	 SIGNAL  rdid_opcode :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  reach_max_cnt :	STD_LOGIC;
	 SIGNAL  read_buf :	STD_LOGIC;
	 SIGNAL  read_bufdly :	STD_LOGIC;
	 SIGNAL  read_data_reg_in_wire :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  read_opcode :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  read_rdid_wire :	STD_LOGIC;
	 SIGNAL  read_sid_wire :	STD_LOGIC;
	 SIGNAL  read_status_wire :	STD_LOGIC;
	 SIGNAL  read_wire :	STD_LOGIC;
	 SIGNAL  rsid_opcode :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  rsid_sdoin :	STD_LOGIC;
	 SIGNAL  rstat_opcode :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  scein_wire :	STD_LOGIC;
	 SIGNAL  sdoin_wire :	STD_LOGIC;
	 SIGNAL  sec_erase_wire :	STD_LOGIC;
	 SIGNAL  sec_protect_wire :	STD_LOGIC;
	 SIGNAL  secprot_opcode :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  secprot_sdoin :	STD_LOGIC;
	 SIGNAL  serase_opcode :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  shift_bytes_wire :	STD_LOGIC;
	 SIGNAL  shift_opcode :	STD_LOGIC;
	 SIGNAL  shift_opdata :	STD_LOGIC;
	 SIGNAL  shift_pgwr_data :	STD_LOGIC;
	 SIGNAL  st_busy_wire :	STD_LOGIC;
	 SIGNAL  stage2_wire :	STD_LOGIC;
	 SIGNAL  stage3_wire :	STD_LOGIC;
	 SIGNAL  stage4_wire :	STD_LOGIC;
	 SIGNAL  start_poll :	STD_LOGIC;
	 SIGNAL  start_sppoll :	STD_LOGIC;
	 SIGNAL  start_wrpoll :	STD_LOGIC;
	 SIGNAL  to_sdoin_wire :	STD_LOGIC;
	 SIGNAL  wren_opcode :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wren_wire :	STD_LOGIC;
	 SIGNAL  write_opcode :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  write_prot_true :	STD_LOGIC;
	 SIGNAL  write_sdoin :	STD_LOGIC;
	 SIGNAL  write_wire :	STD_LOGIC;
	 SIGNAL  wire_w_addr_range279w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_addr_range274w	:	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  wire_w_berase_opcode_range183w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_berase_opcode_range134w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_dataout_wire_range316w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_fast_read_opcode_range191w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_fast_read_opcode_range152w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_pagewr_buf_not_empty_range422w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_pagewr_buf_not_empty_range426w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_pagewr_buf_not_empty_range429w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_pagewr_buf_not_empty_range432w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_pagewr_buf_not_empty_range435w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_pagewr_buf_not_empty_range438w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_pagewr_buf_not_empty_range441w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_pagewr_buf_not_empty_range444w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_pagewr_buf_not_empty_range53w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_rdid_opcode_range197w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_rdid_opcode_range163w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_read_opcode_range193w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_read_opcode_range155w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_rsid_opcode_range199w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_rsid_opcode_range166w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_rstat_opcode_range187w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_rstat_opcode_range144w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_secprot_opcode_range195w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_secprot_opcode_range158w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_serase_opcode_range185w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_serase_opcode_range139w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_wren_opcode_range181w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_wren_opcode_range131w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_write_opcode_range189w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_write_opcode_range147w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 COMPONENT  a_graycounter
	 GENERIC 
	 (
		PVALUE	:	NATURAL := 0;
		WIDTH	:	NATURAL := 8;
		lpm_type	:	STRING := "a_graycounter"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		clk_en	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC;
		cnt_en	:	IN STD_LOGIC := '1';
		q	:	OUT STD_LOGIC_VECTOR(width-1 DOWNTO 0);
		qbin	:	OUT STD_LOGIC_VECTOR(width-1 DOWNTO 0);
		sclr	:	IN STD_LOGIC := '0';
		updown	:	IN STD_LOGIC := '1'
	 ); 
	 END COMPONENT;
	 COMPONENT  lpm_compare
	 GENERIC 
	 (
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_REPRESENTATION	:	STRING := "UNSIGNED";
		LPM_WIDTH	:	NATURAL;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_compare"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		aeb	:	OUT STD_LOGIC;
		agb	:	OUT STD_LOGIC;
		ageb	:	OUT STD_LOGIC;
		alb	:	OUT STD_LOGIC;
		aleb	:	OUT STD_LOGIC;
		aneb	:	OUT STD_LOGIC;
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		dataa	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0')
	 ); 
	 END COMPONENT;
	 COMPONENT  lpm_counter
	 GENERIC 
	 (
		lpm_avalue	:	STRING := "0";
		lpm_direction	:	STRING := "DEFAULT";
		lpm_modulus	:	NATURAL := 0;
		lpm_port_updown	:	STRING := "PORT_CONNECTIVITY";
		lpm_pvalue	:	STRING := "0";
		lpm_svalue	:	STRING := "0";
		lpm_width	:	NATURAL;
		lpm_type	:	STRING := "lpm_counter"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		aload	:	IN STD_LOGIC := '0';
		aset	:	IN STD_LOGIC := '0';
		cin	:	IN STD_LOGIC := '1';
		clk_en	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC;
		cnt_en	:	IN STD_LOGIC := '1';
		cout	:	OUT STD_LOGIC;
		data	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		eq	:	OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
		q	:	OUT STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0);
		sclr	:	IN STD_LOGIC := '0';
		sload	:	IN STD_LOGIC := '0';
		sset	:	IN STD_LOGIC := '0';
		updown	:	IN STD_LOGIC := '1'
	 ); 
	 END COMPONENT;
	 COMPONENT  scfifo
	 GENERIC 
	 (
		ADD_RAM_OUTPUT_REGISTER	:	STRING := "OFF";
		ALLOW_RWCYCLE_WHEN_FULL	:	STRING := "OFF";
		ALMOST_EMPTY_VALUE	:	NATURAL := 0;
		ALMOST_FULL_VALUE	:	NATURAL := 0;
		LPM_NUMWORDS	:	NATURAL;
		LPM_SHOWAHEAD	:	STRING := "OFF";
		LPM_WIDTH	:	NATURAL;
		LPM_WIDTHU	:	NATURAL := 1;
		OVERFLOW_CHECKING	:	STRING := "ON";
		UNDERFLOW_CHECKING	:	STRING := "ON";
		USE_EAB	:	STRING := "ON";
		lpm_type	:	STRING := "scfifo"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		almost_empty	:	OUT STD_LOGIC;
		almost_full	:	OUT STD_LOGIC;
		clock	:	IN STD_LOGIC;
		data	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0);
		empty	:	OUT STD_LOGIC;
		full	:	OUT STD_LOGIC;
		q	:	OUT STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0);
		rdreq	:	IN STD_LOGIC;
		sclr	:	IN STD_LOGIC := '0';
		usedw	:	OUT STD_LOGIC_VECTOR(LPM_WIDTHU-1 DOWNTO 0);
		wrreq	:	IN STD_LOGIC
	 ); 
	 END COMPONENT;
	 COMPONENT  arriaii_asmiblock
	 PORT
	 ( 
		data0in	:	IN STD_LOGIC := '0';
		data0out	:	OUT STD_LOGIC;
		dclkin	:	IN STD_LOGIC;
		dclkout	:	OUT STD_LOGIC;
		oe	:	IN STD_LOGIC := '0';
		scein	:	IN STD_LOGIC;
		sceout	:	OUT STD_LOGIC;
		sdoin	:	IN STD_LOGIC;
		sdoout	:	OUT STD_LOGIC
	 ); 
	 END COMPONENT;
 BEGIN

	wire_w383w(0) <= wire_w_lg_w_lg_w_lg_w_lg_end_operation379w380w381w382w(0) AND wire_w_lg_do_sec_prot375w(0);
	wire_w348w(0) <= wire_w_lg_w_lg_w_lg_w_lg_do_read301w345w346w347w(0) AND end_read_byte;
	wire_w_lg_w_lg_w_lg_w_lg_end_operation379w380w381w382w(0) <= wire_w_lg_w_lg_w_lg_end_operation379w380w381w(0) AND wire_w_lg_do_bulk_erase376w(0);
	wire_w_lg_w_lg_w_lg_w_lg_load_opcode135w136w137w184w(0) <= wire_w_lg_w_lg_w_lg_load_opcode135w136w137w(0) AND wire_w_berase_opcode_range183w(0);
	loop0 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_w_lg_w_lg_load_opcode135w136w137w138w(i) <= wire_w_lg_w_lg_w_lg_load_opcode135w136w137w(0) AND wire_w_berase_opcode_range134w(i);
	END GENERATE loop0;
	wire_w_lg_w_lg_w_lg_w_lg_load_opcode140w141w142w186w(0) <= wire_w_lg_w_lg_w_lg_load_opcode140w141w142w(0) AND wire_w_serase_opcode_range185w(0);
	loop1 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_w_lg_w_lg_load_opcode140w141w142w143w(i) <= wire_w_lg_w_lg_w_lg_load_opcode140w141w142w(0) AND wire_w_serase_opcode_range139w(i);
	END GENERATE loop1;
	wire_w_lg_w_lg_w_lg_w_lg_load_opcode159w160w161w196w(0) <= wire_w_lg_w_lg_w_lg_load_opcode159w160w161w(0) AND wire_w_secprot_opcode_range195w(0);
	loop2 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_w_lg_w_lg_load_opcode159w160w161w162w(i) <= wire_w_lg_w_lg_w_lg_load_opcode159w160w161w(0) AND wire_w_secprot_opcode_range158w(i);
	END GENERATE loop2;
	wire_w_lg_w_lg_w_lg_w_lg_do_read245w246w247w248w(0) <= wire_w_lg_w_lg_w_lg_do_read245w246w247w(0) AND end_one_cycle;
	wire_w_lg_w_lg_w_lg_w_lg_do_write378w552w553w554w(0) <= wire_w_lg_w_lg_w_lg_do_write378w552w553w(0) AND end_operation;
	wire_w555w(0) <= wire_w_lg_w_lg_w_lg_w_lg_do_write57w58w548w549w(0) AND end_operation;
	wire_w_lg_w_lg_w_lg_w_lg_do_read301w345w346w347w(0) <= wire_w_lg_w_lg_w_lg_do_read301w345w346w(0) AND end_one_cyc_pos;
	wire_w_lg_w_lg_w_lg_do_sec_erase289w290w291w(0) <= wire_w_lg_w_lg_do_sec_erase289w290w(0) AND end_operation;
	wire_w_lg_w_lg_w_lg_end_operation379w380w381w(0) <= wire_w_lg_w_lg_end_operation379w380w(0) AND wire_w_lg_do_sec_erase377w(0);
	wire_w_lg_w_lg_w_lg_load_opcode135w136w137w(0) <= wire_w_lg_w_lg_load_opcode135w136w(0) AND wire_w_lg_do_read_stat38w(0);
	wire_w_lg_w_lg_w_lg_load_opcode140w141w142w(0) <= wire_w_lg_w_lg_load_opcode140w141w(0) AND wire_w_lg_do_read_stat38w(0);
	wire_w_lg_w_lg_w_lg_load_opcode159w160w161w(0) <= wire_w_lg_w_lg_load_opcode159w160w(0) AND wire_w_lg_do_read_stat38w(0);
	wire_w_lg_w_lg_w_lg_do_read245w246w247w(0) <= wire_w_lg_w_lg_do_read245w246w(0) AND wire_w_lg_w_lg_do_write48w243w(0);
	wire_w_lg_w_lg_w_lg_do_read245w246w292w(0) <= wire_w_lg_w_lg_do_read245w246w(0) AND clr_write_wire;
	wire_w_lg_w_lg_w_lg_do_write378w552w553w(0) <= wire_w_lg_w_lg_do_write378w552w(0) AND wire_w_lg_do_bulk_erase376w(0);
	wire_w_lg_w_lg_w_lg_w_lg_do_write57w58w548w549w(0) <= wire_w_lg_w_lg_w_lg_do_write57w58w548w(0) AND wire_wrstage_cntr_w_lg_w_q_range460w461w(0);
	wire_w_lg_w_lg_w_lg_do_read301w345w346w(0) <= wire_w_lg_w_lg_do_read301w345w(0) AND wire_stage_cntr_w_lg_w_q_range81w86w(0);
	wire_w_lg_w_lg_bp2_wire477w478w(0) <= wire_w_lg_bp2_wire477w(0) AND bp0_wire;
	wire_w_lg_w_lg_do_polling389w390w(0) <= wire_w_lg_do_polling389w(0) AND stage3_dly_reg;
	wire_w_lg_w_lg_do_sec_erase289w290w(0) <= wire_w_lg_do_sec_erase289w(0) AND wire_w_lg_do_read_stat38w(0);
	wire_w_lg_w_lg_do_write148w149w(0) <= wire_w_lg_do_write148w(0) AND wire_w_lg_do_wren39w(0);
	wire_w_lg_w_lg_do_write48w226w(0) <= wire_w_lg_do_write48w(0) AND end_pgwr_data;
	wire_w_lg_w_lg_end_operation379w380w(0) <= wire_w_lg_end_operation379w(0) AND wire_w_lg_do_write378w(0);
	wire_w_lg_w_lg_load_opcode150w190w(0) <= wire_w_lg_load_opcode150w(0) AND wire_w_write_opcode_range189w(0);
	loop3 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_load_opcode150w151w(i) <= wire_w_lg_load_opcode150w(0) AND wire_w_write_opcode_range147w(i);
	END GENERATE loop3;
	wire_w_lg_w_lg_load_opcode135w136w(0) <= wire_w_lg_load_opcode135w(0) AND wire_w_lg_do_wren39w(0);
	wire_w_lg_w_lg_load_opcode153w192w(0) <= wire_w_lg_load_opcode153w(0) AND wire_w_fast_read_opcode_range191w(0);
	loop4 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_load_opcode153w154w(i) <= wire_w_lg_load_opcode153w(0) AND wire_w_fast_read_opcode_range152w(i);
	END GENERATE loop4;
	wire_w_lg_w_lg_load_opcode156w194w(0) <= wire_w_lg_load_opcode156w(0) AND wire_w_read_opcode_range193w(0);
	loop5 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_load_opcode156w157w(i) <= wire_w_lg_load_opcode156w(0) AND wire_w_read_opcode_range155w(i);
	END GENERATE loop5;
	wire_w_lg_w_lg_load_opcode164w198w(0) <= wire_w_lg_load_opcode164w(0) AND wire_w_rdid_opcode_range197w(0);
	loop6 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_load_opcode164w165w(i) <= wire_w_lg_load_opcode164w(0) AND wire_w_rdid_opcode_range163w(i);
	END GENERATE loop6;
	wire_w_lg_w_lg_load_opcode167w200w(0) <= wire_w_lg_load_opcode167w(0) AND wire_w_rsid_opcode_range199w(0);
	loop7 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_load_opcode167w168w(i) <= wire_w_lg_load_opcode167w(0) AND wire_w_rsid_opcode_range166w(i);
	END GENERATE loop7;
	wire_w_lg_w_lg_load_opcode145w188w(0) <= wire_w_lg_load_opcode145w(0) AND wire_w_rstat_opcode_range187w(0);
	loop8 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_load_opcode145w146w(i) <= wire_w_lg_load_opcode145w(0) AND wire_w_rstat_opcode_range144w(i);
	END GENERATE loop8;
	wire_w_lg_w_lg_load_opcode140w141w(0) <= wire_w_lg_load_opcode140w(0) AND wire_w_lg_do_wren39w(0);
	wire_w_lg_w_lg_load_opcode159w160w(0) <= wire_w_lg_load_opcode159w(0) AND wire_w_lg_do_wren39w(0);
	wire_w_lg_w_lg_load_opcode132w182w(0) <= wire_w_lg_load_opcode132w(0) AND wire_w_wren_opcode_range181w(0);
	loop9 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_load_opcode132w133w(i) <= wire_w_lg_load_opcode132w(0) AND wire_w_wren_opcode_range131w(i);
	END GENERATE loop9;
	wire_w_lg_w_lg_reach_max_cnt453w454w(0) <= wire_w_lg_reach_max_cnt453w(0) AND wren_wire;
	wire_w_lg_w_lg_start_poll231w232w(0) <= wire_w_lg_start_poll231w(0) AND do_polling;
	wire_w_lg_w_lg_do_read245w246w(0) <= wire_w_lg_do_read245w(0) AND wire_w_lg_do_fast_read244w(0);
	wire_w_lg_w_lg_do_write378w552w(0) <= wire_w_lg_do_write378w(0) AND wire_w_lg_do_sec_erase377w(0);
	loop10 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_read_bufdly408w409w(i) <= wire_w_lg_read_bufdly408w(0) AND wire_pgwrbuf_dataout_w_q_range407w(i);
	END GENERATE loop10;
	wire_w_lg_w_lg_w_lg_do_write57w58w457w(0) <= wire_w_lg_w_lg_do_write57w58w(0) AND end_wrstage;
	wire_w_lg_w_lg_w_lg_do_write57w58w59w(0) <= wire_w_lg_w_lg_do_write57w58w(0) AND write_prot_true;
	wire_w_lg_w_lg_w_lg_do_write57w58w548w(0) <= wire_w_lg_w_lg_do_write57w58w(0) AND wire_wrstage_cntr_w_q_range462w(0);
	wire_w_lg_w_lg_do_read301w345w(0) <= wire_w_lg_do_read301w(0) AND wire_stage_cntr_w_q_range82w(0);
	wire_w_lg_w_lg_do_write57w282w(0) <= wire_w_lg_do_write57w(0) AND do_memadd;
	wire_w_lg_w_lg_end_operation391w392w(0) <= wire_w_lg_end_operation391w(0) AND do_read_stat;
	wire_w_lg_w_lg_rden_wire286w287w(0) <= wire_w_lg_rden_wire286w(0) AND not_busy;
	wire_w_lg_bp2_wire477w(0) <= bp2_wire AND bp1_wire;
	wire_w_lg_do_bulk_erase227w(0) <= do_bulk_erase AND wire_w_lg_do_read_stat38w(0);
	wire_w_lg_do_polling389w(0) <= do_polling AND end_one_cyc_pos;
	wire_w_lg_do_sec_erase289w(0) <= do_sec_erase AND wire_w_lg_do_wren39w(0);
	wire_w_lg_do_write148w(0) <= do_write AND wire_w_lg_do_read_stat38w(0);
	wire_w_lg_do_write55w(0) <= do_write AND wire_w_lg_w_pagewr_buf_not_empty_range53w54w(0);
	wire_w_lg_do_write48w(0) <= do_write AND shift_pgwr_data;
	wire_w_lg_end_operation379w(0) <= end_operation AND do_read_stat;
	wire_w_lg_load_opcode150w(0) <= load_opcode AND wire_w_lg_w_lg_do_write148w149w(0);
	wire_w_lg_load_opcode135w(0) <= load_opcode AND do_bulk_erase;
	wire_w_lg_load_opcode153w(0) <= load_opcode AND do_fast_read;
	wire_w_lg_load_opcode156w(0) <= load_opcode AND do_read;
	wire_w_lg_load_opcode164w(0) <= load_opcode AND do_read_rdid;
	wire_w_lg_load_opcode167w(0) <= load_opcode AND do_read_sid;
	wire_w_lg_load_opcode145w(0) <= load_opcode AND do_read_stat;
	wire_w_lg_load_opcode140w(0) <= load_opcode AND do_sec_erase;
	wire_w_lg_load_opcode159w(0) <= load_opcode AND do_sec_prot;
	wire_w_lg_load_opcode132w(0) <= load_opcode AND do_wren;
	wire_w_lg_not_busy280w(0) <= not_busy AND wire_w_addr_range279w(0);
	loop11 : FOR i IN 0 TO 22 GENERATE 
		wire_w_lg_not_busy275w(i) <= not_busy AND wire_w_addr_range274w(i);
	END GENERATE loop11;
	wire_w_lg_reach_max_cnt453w(0) <= reach_max_cnt AND shift_bytes_wire;
	wire_w_lg_read_bufdly416w(0) <= read_bufdly AND wire_scfifo3_w_q_range415w(0);
	loop12 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_read_bufdly411w(i) <= read_bufdly AND wire_scfifo3_w_q_range410w(i);
	END GENERATE loop12;
	loop13 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_shift_opcode130w(i) <= shift_opcode AND wire_asmi_opcode_reg_w_q_range129w(i);
	END GENERATE loop13;
	wire_w_lg_stage3_wire285w(0) <= stage3_wire AND wire_w_lg_w_lg_w_lg_w_lg_do_write57w282w283w284w(0);
	wire_w_lg_stage3_wire312w(0) <= stage3_wire AND wire_w_lg_do_read_stat311w(0);
	loop14 : FOR i IN 0 TO 22 GENERATE 
		wire_w_lg_stage3_wire273w(i) <= stage3_wire AND wire_addr_reg_w_q_range272w(i);
	END GENERATE loop14;
	wire_w_lg_stage4_wire314w(0) <= stage4_wire AND wire_w_lg_w_lg_do_read301w313w(0);
	wire_w_lg_start_poll231w(0) <= start_poll AND do_read_stat;
	wire_w_lg_w_lg_do_write48w243w(0) <= NOT wire_w_lg_do_write48w(0);
	wire_w_lg_bp0_wire479w(0) <= NOT bp0_wire;
	wire_w_lg_bp1_wire483w(0) <= NOT bp1_wire;
	wire_w_lg_bp2_wire494w(0) <= NOT bp2_wire;
	wire_w_lg_buf_empty524w(0) <= NOT buf_empty;
	wire_w_lg_busy_wire1w(0) <= NOT busy_wire;
	wire_w_lg_clkin_wire80w(0) <= NOT clkin_wire;
	wire_w_lg_do_bulk_erase376w(0) <= NOT do_bulk_erase;
	wire_w_lg_do_fast_read244w(0) <= NOT do_fast_read;
	wire_w_lg_do_memadd298w(0) <= NOT do_memadd;
	wire_w_lg_do_polling239w(0) <= NOT do_polling;
	wire_w_lg_do_read245w(0) <= NOT do_read;
	wire_w_lg_do_read_rdid37w(0) <= NOT do_read_rdid;
	wire_w_lg_do_read_stat38w(0) <= NOT do_read_stat;
	wire_w_lg_do_sec_erase377w(0) <= NOT do_sec_erase;
	wire_w_lg_do_sec_prot375w(0) <= NOT do_sec_prot;
	wire_w_lg_do_wren39w(0) <= NOT do_wren;
	wire_w_lg_do_write378w(0) <= NOT do_write;
	wire_w_lg_end_add_cycle67w(0) <= NOT end_add_cycle;
	wire_w_lg_end_fast_read61w(0) <= NOT end_fast_read;
	wire_w_lg_end_ophdly35w(0) <= NOT end_ophdly;
	wire_w_lg_end_pgwr_data47w(0) <= NOT end_pgwr_data;
	wire_w_lg_end_read64w(0) <= NOT end_read;
	wire_w_lg_rden_wire360w(0) <= NOT rden_wire;
	wire_w_lg_reach_max_cnt418w(0) <= NOT reach_max_cnt;
	wire_w_lg_read_bufdly408w(0) <= NOT read_bufdly;
	wire_w_lg_read_rdid_wire10w(0) <= NOT read_rdid_wire;
	wire_w_lg_read_sid_wire9w(0) <= NOT read_sid_wire;
	wire_w_lg_read_status_wire23w(0) <= NOT read_status_wire;
	wire_w_lg_sec_protect_wire8w(0) <= NOT sec_protect_wire;
	wire_w_lg_st_busy_wire95w(0) <= NOT st_busy_wire;
	wire_w_lg_write_prot_true456w(0) <= NOT write_prot_true;
	wire_w_lg_write_wire18w(0) <= NOT write_wire;
	wire_w_lg_w_pagewr_buf_not_empty_range53w54w(0) <= NOT wire_w_pagewr_buf_not_empty_range53w(0);
	wire_w_lg_w555w556w(0) <= wire_w555w(0) OR write_prot_true;
	wire_w_lg_w_lg_w_lg_load_opcode167w200w201w(0) <= wire_w_lg_w_lg_load_opcode167w200w(0) OR wire_w_lg_w_lg_load_opcode164w198w(0);
	loop15 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_w_lg_load_opcode167w168w169w(i) <= wire_w_lg_w_lg_load_opcode167w168w(i) OR wire_w_lg_w_lg_load_opcode164w165w(i);
	END GENERATE loop15;
	wire_w_lg_w_lg_w_lg_do_write57w282w283w(0) <= wire_w_lg_w_lg_do_write57w282w(0) OR do_read;
	wire_w_lg_w_lg_w_lg_rden_wire286w287w288w(0) <= wire_w_lg_w_lg_rden_wire286w287w(0) OR wire_w_lg_stage3_wire285w(0);
	loop16 : FOR i IN 0 TO 22 GENERATE 
		wire_w_lg_w_lg_not_busy275w276w(i) <= wire_w_lg_not_busy275w(i) OR wire_w_lg_stage3_wire273w(i);
	END GENERATE loop16;
	loop17 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_read_bufdly411w412w(i) <= wire_w_lg_read_bufdly411w(i) OR wire_w_lg_w_lg_read_bufdly408w409w(i);
	END GENERATE loop17;
	wire_w_lg_w_lg_stage4_wire314w315w(0) <= wire_w_lg_stage4_wire314w(0) OR wire_w_lg_stage3_wire312w(0);
	wire_w_lg_w_lg_w_lg_w_lg_load_opcode167w200w201w202w(0) <= wire_w_lg_w_lg_w_lg_load_opcode167w200w201w(0) OR wire_w_lg_w_lg_w_lg_w_lg_load_opcode159w160w161w196w(0);
	loop18 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_w_lg_w_lg_load_opcode167w168w169w170w(i) <= wire_w_lg_w_lg_w_lg_load_opcode167w168w169w(i) OR wire_w_lg_w_lg_w_lg_w_lg_load_opcode159w160w161w162w(i);
	END GENERATE loop18;
	wire_w_lg_w_lg_w_lg_w_lg_do_write57w282w283w284w(0) <= wire_w_lg_w_lg_w_lg_do_write57w282w283w(0) OR do_fast_read;
	wire_w203w(0) <= wire_w_lg_w_lg_w_lg_w_lg_load_opcode167w200w201w202w(0) OR wire_w_lg_w_lg_load_opcode156w194w(0);
	loop19 : FOR i IN 0 TO 6 GENERATE 
		wire_w171w(i) <= wire_w_lg_w_lg_w_lg_w_lg_load_opcode167w168w169w170w(i) OR wire_w_lg_w_lg_load_opcode156w157w(i);
	END GENERATE loop19;
	wire_w_lg_w203w204w(0) <= wire_w203w(0) OR wire_w_lg_w_lg_load_opcode153w192w(0);
	loop20 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w171w172w(i) <= wire_w171w(i) OR wire_w_lg_w_lg_load_opcode153w154w(i);
	END GENERATE loop20;
	wire_w_lg_w_lg_w203w204w205w(0) <= wire_w_lg_w203w204w(0) OR wire_w_lg_w_lg_load_opcode150w190w(0);
	loop21 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_w171w172w173w(i) <= wire_w_lg_w171w172w(i) OR wire_w_lg_w_lg_load_opcode150w151w(i);
	END GENERATE loop21;
	wire_w_lg_w_lg_w_lg_w203w204w205w206w(0) <= wire_w_lg_w_lg_w203w204w205w(0) OR wire_w_lg_w_lg_load_opcode145w188w(0);
	loop22 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_w_lg_w171w172w173w174w(i) <= wire_w_lg_w_lg_w171w172w173w(i) OR wire_w_lg_w_lg_load_opcode145w146w(i);
	END GENERATE loop22;
	wire_w_lg_w_lg_w_lg_w_lg_w203w204w205w206w207w(0) <= wire_w_lg_w_lg_w_lg_w203w204w205w206w(0) OR wire_w_lg_w_lg_w_lg_w_lg_load_opcode140w141w142w186w(0);
	loop23 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_w_lg_w_lg_w171w172w173w174w175w(i) <= wire_w_lg_w_lg_w_lg_w171w172w173w174w(i) OR wire_w_lg_w_lg_w_lg_w_lg_load_opcode140w141w142w143w(i);
	END GENERATE loop23;
	wire_w_lg_w_lg_w_lg_w_lg_w_lg_w203w204w205w206w207w208w(0) <= wire_w_lg_w_lg_w_lg_w_lg_w203w204w205w206w207w(0) OR wire_w_lg_w_lg_w_lg_w_lg_load_opcode135w136w137w184w(0);
	loop24 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_w_lg_w_lg_w_lg_w171w172w173w174w175w176w(i) <= wire_w_lg_w_lg_w_lg_w_lg_w171w172w173w174w175w(i) OR wire_w_lg_w_lg_w_lg_w_lg_load_opcode135w136w137w138w(i);
	END GENERATE loop24;
	wire_w209w(0) <= wire_w_lg_w_lg_w_lg_w_lg_w_lg_w203w204w205w206w207w208w(0) OR wire_w_lg_w_lg_load_opcode132w182w(0);
	loop25 : FOR i IN 0 TO 6 GENERATE 
		wire_w177w(i) <= wire_w_lg_w_lg_w_lg_w_lg_w_lg_w171w172w173w174w175w176w(i) OR wire_w_lg_w_lg_load_opcode132w133w(i);
	END GENERATE loop25;
	loop26 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w177w178w(i) <= wire_w177w(i) OR wire_w_lg_shift_opcode130w(i);
	END GENERATE loop26;
	wire_w117w(0) <= wire_w_lg_w_lg_w_lg_w_lg_do_read_sid113w114w115w116w(0) OR do_read_rdid;
	wire_w_lg_w_lg_w_lg_w_lg_do_read_sid113w114w115w116w(0) <= wire_w_lg_w_lg_w_lg_do_read_sid113w114w115w(0) OR do_sec_erase;
	wire_w_lg_w_lg_w_lg_do_read301w302w303w(0) <= wire_w_lg_w_lg_do_read301w302w(0) OR do_sec_erase;
	wire_w_lg_w_lg_w_lg_do_read_sid113w114w115w(0) <= wire_w_lg_w_lg_do_read_sid113w114w(0) OR do_write;
	wire_w_lg_w_lg_do_read301w313w(0) <= wire_w_lg_do_read301w(0) OR do_read_sid;
	wire_w_lg_w_lg_do_read301w302w(0) <= wire_w_lg_do_read301w(0) OR do_write;
	wire_w_lg_w_lg_do_read_sid113w114w(0) <= wire_w_lg_do_read_sid113w(0) OR do_fast_read;
	wire_w_lg_w_lg_do_sec_erase468w469w(0) <= wire_w_lg_do_sec_erase468w(0) OR do_bulk_erase;
	wire_w_lg_w_lg_do_write57w58w(0) <= wire_w_lg_do_write57w(0) OR do_bulk_erase;
	wire_w_lg_data0out_wire317w(0) <= data0out_wire OR wire_w_dataout_wire_range316w(0);
	wire_w_lg_do_read301w(0) <= do_read OR do_fast_read;
	wire_w_lg_do_read_sid113w(0) <= do_read_sid OR do_read;
	wire_w_lg_do_read_stat311w(0) <= do_read_stat OR do_read_rdid;
	wire_w_lg_do_sec_erase468w(0) <= do_sec_erase OR do_write;
	wire_w_lg_do_wren228w(0) <= do_wren OR wire_w_lg_do_bulk_erase227w(0);
	wire_w_lg_do_write57w(0) <= do_write OR do_sec_erase;
	wire_w_lg_end_operation391w(0) <= end_operation OR wire_w_lg_w_lg_do_polling389w390w(0);
	wire_w_lg_load_opcode211w(0) <= load_opcode OR shift_opcode;
	wire_w_lg_rden_wire286w(0) <= rden_wire OR wren_wire;
	wire_w_lg_read_bufdly406w(0) <= read_bufdly OR shift_pgwr_data;
	wire_w_lg_w_pagewr_buf_not_empty_range422w425w(0) <= wire_w_pagewr_buf_not_empty_range422w(0) OR wire_pgwr_data_cntr_w_q_range424w(0);
	wire_w_lg_w_pagewr_buf_not_empty_range426w428w(0) <= wire_w_pagewr_buf_not_empty_range426w(0) OR wire_pgwr_data_cntr_w_q_range427w(0);
	wire_w_lg_w_pagewr_buf_not_empty_range429w431w(0) <= wire_w_pagewr_buf_not_empty_range429w(0) OR wire_pgwr_data_cntr_w_q_range430w(0);
	wire_w_lg_w_pagewr_buf_not_empty_range432w434w(0) <= wire_w_pagewr_buf_not_empty_range432w(0) OR wire_pgwr_data_cntr_w_q_range433w(0);
	wire_w_lg_w_pagewr_buf_not_empty_range435w437w(0) <= wire_w_pagewr_buf_not_empty_range435w(0) OR wire_pgwr_data_cntr_w_q_range436w(0);
	wire_w_lg_w_pagewr_buf_not_empty_range438w440w(0) <= wire_w_pagewr_buf_not_empty_range438w(0) OR wire_pgwr_data_cntr_w_q_range439w(0);
	wire_w_lg_w_pagewr_buf_not_empty_range441w443w(0) <= wire_w_pagewr_buf_not_empty_range441w(0) OR wire_pgwr_data_cntr_w_q_range442w(0);
	wire_w_lg_w_pagewr_buf_not_empty_range444w446w(0) <= wire_w_pagewr_buf_not_empty_range444w(0) OR wire_pgwr_data_cntr_w_q_range445w(0);
	be_write_prot <= (do_bulk_erase AND (((bp3_wire OR bp2_wire) OR bp1_wire) OR bp0_wire));
	berase_opcode <= (OTHERS => '0');
	bp0_wire <= statreg_int(2);
	bp1_wire <= statreg_int(3);
	bp2_wire <= statreg_int(4);
	bp3_wire <= statreg_int(6);
	buf_empty <= buf_empty_reg;
	busy <= busy_wire;
	busy_wire <= ((((((((do_read_rdid OR do_read_sid) OR do_read) OR do_fast_read) OR do_write) OR do_sec_prot) OR do_read_stat) OR do_sec_erase) OR do_bulk_erase);
	clkin_wire <= clkin;
	clr_rdid_wire <= clr_rdid_reg2;
	clr_read_wire <= clr_read_reg2;
	clr_rstat_wire <= clr_rstat_reg2;
	clr_write_wire <= clr_write_reg2;
	cnt_bfend_wire_in <= (wire_gen_cntr_w_lg_w_q_range92w93w(0) AND wire_gen_cntr_q(0));
	data0out_wire <= wire_stratixii_asmiblock2_data0out;
	data_valid <= data_valid_wire;
	data_valid_wire <= dvalid_reg2;
	dataout <= ( read_data_reg(7 DOWNTO 0));
	dataout_wire <= ( "0000");
	do_bulk_erase <= '0';
	do_fast_read <= '0';
	do_memadd <= do_wrmemadd_reg;
	do_polling <= (do_write_polling OR do_sprot_polling);
	do_read <= (((wire_w_lg_read_rdid_wire10w(0) AND wire_w_lg_read_sid_wire9w(0)) AND wire_w_lg_sec_protect_wire8w(0)) AND read_wire);
	do_read_rdid <= read_rdid_wire;
	do_read_sid <= '0';
	do_read_stat <= (((((((wire_w_lg_read_rdid_wire10w(0) AND wire_w_lg_read_sid_wire9w(0)) AND wire_w_lg_sec_protect_wire8w(0)) AND (NOT (read_wire OR fast_read_wire))) AND wire_w_lg_write_wire18w(0)) AND read_status_wire) OR do_write_rstat) OR do_sprot_rstat);
	do_sec_erase <= ((((((wire_w_lg_read_rdid_wire10w(0) AND wire_w_lg_read_sid_wire9w(0)) AND wire_w_lg_sec_protect_wire8w(0)) AND (NOT (read_wire OR fast_read_wire))) AND wire_w_lg_write_wire18w(0)) AND wire_w_lg_read_status_wire23w(0)) AND sec_erase_wire);
	do_sec_prot <= '0';
	do_secprot_wren <= '0';
	do_sprot_polling <= '0';
	do_sprot_rstat <= '0';
	do_wren <= (do_write_wren OR do_secprot_wren);
	do_write <= ((((wire_w_lg_read_rdid_wire10w(0) AND wire_w_lg_read_sid_wire9w(0)) AND wire_w_lg_sec_protect_wire8w(0)) AND (NOT (read_wire OR fast_read_wire))) AND write_wire);
	do_write_polling <= wire_w_lg_w_lg_w_lg_w_lg_do_write57w58w548w549w(0);
	do_write_rstat <= write_rstat_reg;
	do_write_wren <= ((NOT wire_wrstage_cntr_q(1)) AND wire_wrstage_cntr_q(0));
	dummy_read_buf <= maxcnt_shift_reg2;
	end1_cyc_gen_cntr_wire <= (wire_gen_cntr_w_lg_w_q_range92w93w(0) AND (NOT wire_gen_cntr_q(0)));
	end1_cyc_normal_in_wire <= (((((((((wire_stage_cntr_w_lg_w_lg_w_q_range81w86w100w(0) AND (NOT wire_gen_cntr_q(2))) AND wire_gen_cntr_q(1)) AND wire_gen_cntr_q(0)) OR wire_stage_cntr_w_lg_w_lg_w_lg_w_lg_w_q_range81w86w100w101w102w(0)) OR (do_read AND end_read)) OR (do_fast_read AND end_fast_read)) OR wire_w_lg_w_lg_w_lg_do_write57w58w59w(0)) OR wire_w_lg_do_write55w(0)) OR ((do_read_stat AND start_poll) AND wire_w_lg_st_busy_wire95w(0)));
	end1_cyc_reg_in_wire <= end1_cyc_normal_in_wire;
	end_add_cycle <= wire_mux211_dataout;
	end_add_cycle_mux_datab_wire <= wire_addbyte_cntr_q(2);
	end_fast_read <= end_read_reg;
	end_one_cyc_pos <= end1_cyc_reg2;
	end_one_cycle <= end1_cyc_reg;
	end_operation <= end_op_reg;
	end_ophdly <= end_op_hdlyreg;
	end_pgwr_data <= end_pgwrop_reg;
	end_read <= end_read_reg;
	end_read_byte <= end_rbyte_reg;
	end_wrstage <= end_operation;
	fast_read_opcode <= (OTHERS => '0');
	fast_read_wire <= '0';
	ill_erase_wire <= ill_erase_reg;
	ill_write_wire <= ill_write_reg;
	illegal_erase <= ill_erase_wire;
	illegal_erase_b4out_wire <= ((do_sec_erase OR do_bulk_erase) AND write_prot_true);
	illegal_write <= ill_write_wire;
	illegal_write_b4out_wire <= ((do_write AND write_prot_true) OR wire_w_lg_do_write55w(0));
	in_operation <= busy_wire;
	load_opcode <= ((((wire_stage_cntr_w_lg_w_q_range82w83w(0) AND wire_stage_cntr_w_lg_w_q_range81w86w(0)) AND (NOT wire_gen_cntr_q(2))) AND wire_gen_cntr_w_lg_w_q_range90w91w(0)) AND wire_gen_cntr_q(0));
	memadd_sdoin <= add_msb_reg;
	not_busy <= busy_det_reg;
	oe_wire <= '0';
	page_size_wire <= "100000000";
	pagewr_buf_not_empty <= ( wire_w_lg_w_pagewr_buf_not_empty_range444w446w & wire_w_lg_w_pagewr_buf_not_empty_range441w443w & wire_w_lg_w_pagewr_buf_not_empty_range438w440w & wire_w_lg_w_pagewr_buf_not_empty_range435w437w & wire_w_lg_w_pagewr_buf_not_empty_range432w434w & wire_w_lg_w_pagewr_buf_not_empty_range429w431w & wire_w_lg_w_pagewr_buf_not_empty_range426w428w & wire_w_lg_w_pagewr_buf_not_empty_range422w425w & wire_pgwr_data_cntr_q(0));
	rden_wire <= rden;
	rdid_load <= (end_operation AND do_read_rdid);
	rdid_opcode <= "10011111";
	rdid_out <= ( rdid_out_reg(7 DOWNTO 0));
	reach_max_cnt <= max_cnt_reg;
	read_buf <= (((((end_one_cycle AND do_write) AND wire_w_lg_do_read_stat38w(0)) AND wire_w_lg_do_wren39w(0)) AND (wire_stage_cntr_w_lg_w_q_range82w87w(0) OR wire_addbyte_cntr_w_lg_w_q_range123w124w(0))) AND wire_w_lg_buf_empty524w(0));
	read_bufdly <= read_bufdly_reg;
	read_data_reg_in_wire <= ( read_dout_reg(7 DOWNTO 0));
	read_opcode <= "00000011";
	read_rdid_wire <= read_rdid_reg;
	read_sid_wire <= '0';
	read_status_wire <= read_status_reg;
	read_wire <= read_reg;
	rsid_opcode <= (OTHERS => '0');
	rsid_sdoin <= '0';
	rstat_opcode <= "00000101";
	scein_wire <= wire_ncs_reg_w_lg_q262w(0);
	sdoin_wire <= to_sdoin_wire;
	sec_erase_wire <= sec_erase_reg;
	sec_protect_wire <= '0';
	secprot_opcode <= (OTHERS => '0');
	secprot_sdoin <= '0';
	serase_opcode <= "11011000";
	shift_bytes_wire <= shift_bytes;
	shift_opcode <= shift_op_reg;
	shift_opdata <= stage2_wire;
	shift_pgwr_data <= shftpgwr_data_reg;
	st_busy_wire <= statreg_int(0);
	stage2_wire <= stage2_reg;
	stage3_wire <= stage3_reg;
	stage4_wire <= stage4_reg;
	start_poll <= (start_wrpoll OR start_sppoll);
	start_sppoll <= '0';
	start_wrpoll <= start_wrpoll_reg2;
	status_out <= ( statreg_out(7 DOWNTO 0));
	to_sdoin_wire <= (((((shift_opdata AND asmi_opcode_reg(7)) OR rsid_sdoin) OR memadd_sdoin) OR write_sdoin) OR secprot_sdoin);
	wren_opcode <= "00000110";
	wren_wire <= wren;
	write_opcode <= "00000010";
	write_prot_true <= write_prot_reg;
	write_sdoin <= ((((do_write AND stage4_wire) AND wire_wrstage_cntr_q(1)) AND wire_wrstage_cntr_q(0)) AND pgwrbuf_dataout(7));
	write_wire <= write_reg;
	wire_w_addr_range279w(0) <= addr(0);
	wire_w_addr_range274w <= addr(23 DOWNTO 1);
	wire_w_berase_opcode_range183w(0) <= berase_opcode(0);
	wire_w_berase_opcode_range134w <= berase_opcode(7 DOWNTO 1);
	wire_w_dataout_wire_range316w(0) <= dataout_wire(1);
	wire_w_fast_read_opcode_range191w(0) <= fast_read_opcode(0);
	wire_w_fast_read_opcode_range152w <= fast_read_opcode(7 DOWNTO 1);
	wire_w_pagewr_buf_not_empty_range422w(0) <= pagewr_buf_not_empty(0);
	wire_w_pagewr_buf_not_empty_range426w(0) <= pagewr_buf_not_empty(1);
	wire_w_pagewr_buf_not_empty_range429w(0) <= pagewr_buf_not_empty(2);
	wire_w_pagewr_buf_not_empty_range432w(0) <= pagewr_buf_not_empty(3);
	wire_w_pagewr_buf_not_empty_range435w(0) <= pagewr_buf_not_empty(4);
	wire_w_pagewr_buf_not_empty_range438w(0) <= pagewr_buf_not_empty(5);
	wire_w_pagewr_buf_not_empty_range441w(0) <= pagewr_buf_not_empty(6);
	wire_w_pagewr_buf_not_empty_range444w(0) <= pagewr_buf_not_empty(7);
	wire_w_pagewr_buf_not_empty_range53w(0) <= pagewr_buf_not_empty(8);
	wire_w_rdid_opcode_range197w(0) <= rdid_opcode(0);
	wire_w_rdid_opcode_range163w <= rdid_opcode(7 DOWNTO 1);
	wire_w_read_opcode_range193w(0) <= read_opcode(0);
	wire_w_read_opcode_range155w <= read_opcode(7 DOWNTO 1);
	wire_w_rsid_opcode_range199w(0) <= rsid_opcode(0);
	wire_w_rsid_opcode_range166w <= rsid_opcode(7 DOWNTO 1);
	wire_w_rstat_opcode_range187w(0) <= rstat_opcode(0);
	wire_w_rstat_opcode_range144w <= rstat_opcode(7 DOWNTO 1);
	wire_w_secprot_opcode_range195w(0) <= secprot_opcode(0);
	wire_w_secprot_opcode_range158w <= secprot_opcode(7 DOWNTO 1);
	wire_w_serase_opcode_range185w(0) <= serase_opcode(0);
	wire_w_serase_opcode_range139w <= serase_opcode(7 DOWNTO 1);
	wire_w_wren_opcode_range181w(0) <= wren_opcode(0);
	wire_w_wren_opcode_range131w <= wren_opcode(7 DOWNTO 1);
	wire_w_write_opcode_range189w(0) <= write_opcode(0);
	wire_w_write_opcode_range147w <= write_opcode(7 DOWNTO 1);
	wire_addbyte_cntr_w_lg_w_q_range123w124w(0) <= wire_addbyte_cntr_w_q_range123w(0) AND wire_addbyte_cntr_w_lg_w_q_range121w122w(0);
	wire_addbyte_cntr_w_lg_w_q_range121w122w(0) <= NOT wire_addbyte_cntr_w_q_range121w(0);
	wire_addbyte_cntr_clk_en <= wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range82w85w118w119w(0);
	wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range82w85w118w119w(0) <= wire_stage_cntr_w_lg_w_lg_w_q_range82w85w118w(0) AND wire_w117w(0);
	wire_addbyte_cntr_clock <= wire_w_lg_clkin_wire80w(0);
	wire_addbyte_cntr_w_q_range121w(0) <= wire_addbyte_cntr_q(0);
	wire_addbyte_cntr_w_q_range123w(0) <= wire_addbyte_cntr_q(1);
	addbyte_cntr :  a_graycounter
	  GENERIC MAP (
		WIDTH => 3
	  )
	  PORT MAP ( 
		aclr => end_operation,
		clk_en => wire_addbyte_cntr_clk_en,
		clock => wire_addbyte_cntr_clock,
		q => wire_addbyte_cntr_q
	  );
	wire_gen_cntr_w_lg_w_q_range92w93w(0) <= wire_gen_cntr_w_q_range92w(0) AND wire_gen_cntr_w_lg_w_q_range90w91w(0);
	wire_gen_cntr_w_lg_w_q_range90w91w(0) <= NOT wire_gen_cntr_w_q_range90w(0);
	wire_gen_cntr_clk_en <= wire_w_lg_in_operation36w(0);
	wire_w_lg_in_operation36w(0) <= in_operation AND wire_w_lg_end_ophdly35w(0);
	wire_gen_cntr_w_q_range90w(0) <= wire_gen_cntr_q(1);
	wire_gen_cntr_w_q_range92w(0) <= wire_gen_cntr_q(2);
	gen_cntr :  a_graycounter
	  GENERIC MAP (
		WIDTH => 3
	  )
	  PORT MAP ( 
		aclr => end_one_cycle,
		clk_en => wire_gen_cntr_clk_en,
		clock => clkin_wire,
		q => wire_gen_cntr_q
	  );
	wire_stage_cntr_w_lg_w220w221w(0) <= wire_stage_cntr_w220w(0) AND end_one_cycle;
	wire_stage_cntr_w220w(0) <= wire_stage_cntr_w_lg_w_lg_w_lg_w_lg_w_q_range82w85w217w218w219w(0) AND end_add_cycle;
	wire_stage_cntr_w225w(0) <= wire_stage_cntr_w_lg_w_lg_w_lg_w_lg_w_q_range82w85w222w223w224w(0) AND end_one_cycle;
	wire_stage_cntr_w_lg_w_lg_w_lg_w_lg_w_q_range82w85w217w218w219w(0) <= wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range82w85w217w218w(0) AND wire_w_lg_do_read_stat38w(0);
	wire_stage_cntr_w_lg_w_lg_w_lg_w_lg_w_q_range82w85w222w223w224w(0) <= wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range82w85w222w223w(0) AND wire_w_lg_do_read_stat38w(0);
	wire_stage_cntr_w_lg_w_lg_w_lg_w_lg_w_q_range82w83w84w229w230w(0) <= wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range82w83w84w229w(0) AND end_one_cycle;
	wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range82w87w293w294w(0) <= wire_stage_cntr_w_lg_w_lg_w_q_range82w87w293w(0) AND end_one_cyc_pos;
	wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range82w85w234w235w(0) <= wire_stage_cntr_w_lg_w_lg_w_q_range82w85w234w(0) AND end_one_cycle;
	wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range82w85w240w241w(0) <= wire_stage_cntr_w_lg_w_lg_w_q_range82w85w240w(0) AND end_one_cycle;
	wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range82w85w217w218w(0) <= wire_stage_cntr_w_lg_w_lg_w_q_range82w85w217w(0) AND wire_w_lg_do_wren39w(0);
	wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range82w85w222w223w(0) <= wire_stage_cntr_w_lg_w_lg_w_q_range82w85w222w(0) AND wire_w_lg_do_wren39w(0);
	wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range82w83w84w229w(0) <= wire_stage_cntr_w_lg_w_lg_w_q_range82w83w84w(0) AND wire_w_lg_do_wren228w(0);
	wire_stage_cntr_w_lg_w_lg_w_q_range82w87w293w(0) <= wire_stage_cntr_w_lg_w_q_range82w87w(0) AND end_add_cycle;
	wire_stage_cntr_w_lg_w_lg_w_q_range82w85w234w(0) <= wire_stage_cntr_w_lg_w_q_range82w85w(0) AND do_read_rdid;
	wire_stage_cntr_w_lg_w_lg_w_q_range82w85w240w(0) <= wire_stage_cntr_w_lg_w_q_range82w85w(0) AND do_read_stat;
	wire_stage_cntr_w_lg_w_lg_w_q_range82w85w217w(0) <= wire_stage_cntr_w_lg_w_q_range82w85w(0) AND do_sec_erase;
	wire_stage_cntr_w_lg_w_lg_w_q_range82w85w222w(0) <= wire_stage_cntr_w_lg_w_q_range82w85w(0) AND do_sec_prot;
	wire_stage_cntr_w_lg_w_lg_w_q_range82w85w118w(0) <= wire_stage_cntr_w_lg_w_q_range82w85w(0) AND end_one_cyc_pos;
	wire_stage_cntr_w_lg_w_lg_w_lg_w_lg_w_q_range81w86w100w101w102w(0) <= wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range81w86w100w101w(0) AND end1_cyc_gen_cntr_wire;
	wire_stage_cntr_w_lg_w_lg_w_q_range81w86w100w(0) <= wire_stage_cntr_w_lg_w_q_range81w86w(0) AND wire_stage_cntr_w_lg_w_q_range82w83w(0);
	wire_stage_cntr_w_lg_w_lg_w_q_range82w83w84w(0) <= wire_stage_cntr_w_lg_w_q_range82w83w(0) AND wire_stage_cntr_w_q_range81w(0);
	wire_stage_cntr_w_lg_w_q_range82w87w(0) <= wire_stage_cntr_w_q_range82w(0) AND wire_stage_cntr_w_lg_w_q_range81w86w(0);
	wire_stage_cntr_w_lg_w_q_range82w85w(0) <= wire_stage_cntr_w_q_range82w(0) AND wire_stage_cntr_w_q_range81w(0);
	wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range81w86w100w101w(0) <= NOT wire_stage_cntr_w_lg_w_lg_w_q_range81w86w100w(0);
	wire_stage_cntr_w_lg_w_q_range81w86w(0) <= NOT wire_stage_cntr_w_q_range81w(0);
	wire_stage_cntr_w_lg_w_q_range82w83w(0) <= NOT wire_stage_cntr_w_q_range82w(0);
	wire_stage_cntr_clk_en <= wire_w_lg_w_lg_w_lg_w_lg_w_lg_w74w75w76w77w78w79w(0);
	wire_w_lg_w_lg_w_lg_w_lg_w_lg_w74w75w76w77w78w79w(0) <= (((((((((in_operation AND end_one_cycle) AND (NOT (stage3_wire AND wire_w_lg_end_add_cycle67w(0)))) AND (NOT (stage4_wire AND wire_w_lg_end_read64w(0)))) AND (NOT (stage4_wire AND wire_w_lg_end_fast_read61w(0)))) AND (NOT wire_w_lg_w_lg_w_lg_do_write57w58w59w(0))) AND (NOT wire_w_lg_do_write55w(0))) AND (NOT (stage3_wire AND st_busy_wire))) AND (NOT (wire_w_lg_do_write48w(0) AND wire_w_lg_end_pgwr_data47w(0)))) AND (NOT (stage2_wire AND do_wren))) AND (NOT ((((stage3_wire AND do_sec_erase) AND wire_w_lg_do_wren39w(0)) AND wire_w_lg_do_read_stat38w(0)) AND wire_w_lg_do_read_rdid37w(0)));
	wire_stage_cntr_w_q_range81w(0) <= wire_stage_cntr_q(0);
	wire_stage_cntr_w_q_range82w(0) <= wire_stage_cntr_q(1);
	stage_cntr :  a_graycounter
	  GENERIC MAP (
		WIDTH => 2
	  )
	  PORT MAP ( 
		aclr => end_ophdly,
		clk_en => wire_stage_cntr_clk_en,
		clock => clkin_wire,
		q => wire_stage_cntr_q
	  );
	wire_wrstage_cntr_w_lg_w_q_range462w463w(0) <= wire_wrstage_cntr_w_q_range462w(0) AND wire_wrstage_cntr_w_lg_w_q_range460w461w(0);
	wire_wrstage_cntr_w_lg_w_q_range460w461w(0) <= NOT wire_wrstage_cntr_w_q_range460w(0);
	wire_wrstage_cntr_clk_en <= wire_w459w(0);
	wire_w459w(0) <= (wire_w_lg_w_lg_w_lg_do_write57w58w457w(0) AND wire_w_lg_write_prot_true456w(0)) AND wire_w_lg_st_busy_wire95w(0);
	wire_wrstage_cntr_clock <= wire_w_lg_clkin_wire80w(0);
	wire_wrstage_cntr_w_q_range460w(0) <= wire_wrstage_cntr_q(0);
	wire_wrstage_cntr_w_q_range462w(0) <= wire_wrstage_cntr_q(1);
	wrstage_cntr :  a_graycounter
	  GENERIC MAP (
		WIDTH => 2
	  )
	  PORT MAP ( 
		aclr => clr_write_wire,
		clk_en => wire_wrstage_cntr_clk_en,
		clock => wire_wrstage_cntr_clock,
		q => wire_wrstage_cntr_q
	  );
	PROCESS (clkin_wire, clr_addmsb_reg)
	BEGIN
		IF (clr_addmsb_reg = '1') THEN add_msb_reg <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_add_msb_reg_ena = '1') THEN add_msb_reg <= wire_addr_reg_w_q_range297w(0);
			END IF;
		END IF;
	END PROCESS;
	wire_add_msb_reg_ena <= (((wire_w_lg_w_lg_w_lg_do_read301w302w303w(0) AND (NOT (wire_w_lg_do_write57w(0) AND wire_w_lg_do_memadd298w(0)))) AND wire_stage_cntr_q(1)) AND wire_stage_cntr_q(0));
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(0) = '1') THEN addr_reg(0) <= wire_addr_reg_d(0);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(1) = '1') THEN addr_reg(1) <= wire_addr_reg_d(1);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(2) = '1') THEN addr_reg(2) <= wire_addr_reg_d(2);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(3) = '1') THEN addr_reg(3) <= wire_addr_reg_d(3);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(4) = '1') THEN addr_reg(4) <= wire_addr_reg_d(4);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(5) = '1') THEN addr_reg(5) <= wire_addr_reg_d(5);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(6) = '1') THEN addr_reg(6) <= wire_addr_reg_d(6);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(7) = '1') THEN addr_reg(7) <= wire_addr_reg_d(7);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(8) = '1') THEN addr_reg(8) <= wire_addr_reg_d(8);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(9) = '1') THEN addr_reg(9) <= wire_addr_reg_d(9);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(10) = '1') THEN addr_reg(10) <= wire_addr_reg_d(10);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(11) = '1') THEN addr_reg(11) <= wire_addr_reg_d(11);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(12) = '1') THEN addr_reg(12) <= wire_addr_reg_d(12);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(13) = '1') THEN addr_reg(13) <= wire_addr_reg_d(13);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(14) = '1') THEN addr_reg(14) <= wire_addr_reg_d(14);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(15) = '1') THEN addr_reg(15) <= wire_addr_reg_d(15);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(16) = '1') THEN addr_reg(16) <= wire_addr_reg_d(16);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(17) = '1') THEN addr_reg(17) <= wire_addr_reg_d(17);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(18) = '1') THEN addr_reg(18) <= wire_addr_reg_d(18);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(19) = '1') THEN addr_reg(19) <= wire_addr_reg_d(19);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(20) = '1') THEN addr_reg(20) <= wire_addr_reg_d(20);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(21) = '1') THEN addr_reg(21) <= wire_addr_reg_d(21);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(22) = '1') THEN addr_reg(22) <= wire_addr_reg_d(22);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(23) = '1') THEN addr_reg(23) <= wire_addr_reg_d(23);
			END IF;
		END IF;
	END PROCESS;
	wire_addr_reg_d <= ( wire_w_lg_w_lg_not_busy275w276w & wire_w_lg_not_busy280w);
	loop27 : FOR i IN 0 TO 23 GENERATE
		wire_addr_reg_ena(i) <= wire_w_lg_w_lg_w_lg_rden_wire286w287w288w(0);
	END GENERATE loop27;
	wire_addr_reg_w_lg_w_lg_w_lg_w506w507w508w509w(0) <= wire_addr_reg_w_lg_w_lg_w506w507w508w(0) AND bp0_wire;
	wire_addr_reg_w_lg_w_lg_w506w507w508w(0) <= wire_addr_reg_w_lg_w506w507w(0) AND wire_w_lg_bp1_wire483w(0);
	wire_addr_reg_w_lg_w498w499w(0) <= wire_addr_reg_w498w(0) AND bp0_wire;
	wire_addr_reg_w_lg_w502w503w(0) <= wire_addr_reg_w502w(0) AND bp1_wire;
	wire_addr_reg_w_lg_w506w507w(0) <= wire_addr_reg_w506w(0) AND wire_w_lg_bp2_wire494w(0);
	wire_addr_reg_w498w(0) <= wire_addr_reg_w_lg_w_lg_w_lg_w_lg_w_q_range297w485w490w496w497w(0) AND bp1_wire;
	wire_addr_reg_w502w(0) <= wire_addr_reg_w_lg_w_lg_w_lg_w_lg_w_q_range297w485w490w496w501w(0) AND wire_w_lg_bp2_wire494w(0);
	wire_addr_reg_w506w(0) <= wire_addr_reg_w_lg_w_lg_w_lg_w_lg_w_q_range297w485w490w496w501w(0) AND wire_addr_reg_w_q_range505w(0);
	wire_addr_reg_w_lg_w_lg_w_lg_w_lg_w_q_range297w485w486w487w488w(0) <= wire_addr_reg_w_lg_w_lg_w_lg_w_q_range297w485w486w487w(0) AND bp0_wire;
	wire_addr_reg_w_lg_w_lg_w_lg_w_lg_w_q_range297w485w490w496w497w(0) <= wire_addr_reg_w_lg_w_lg_w_lg_w_q_range297w485w490w496w(0) AND wire_w_lg_bp2_wire494w(0);
	wire_addr_reg_w_lg_w_lg_w_lg_w_lg_w_q_range297w485w490w496w501w(0) <= wire_addr_reg_w_lg_w_lg_w_lg_w_q_range297w485w490w496w(0) AND wire_addr_reg_w_q_range500w(0);
	wire_addr_reg_w_lg_w_lg_w_lg_w_q_range297w485w486w487w(0) <= wire_addr_reg_w_lg_w_lg_w_q_range297w485w486w(0) AND wire_w_lg_bp1_wire483w(0);
	wire_addr_reg_w_lg_w_lg_w_lg_w_q_range297w485w490w491w(0) <= wire_addr_reg_w_lg_w_lg_w_q_range297w485w490w(0) AND bp2_wire;
	wire_addr_reg_w_lg_w_lg_w_lg_w_q_range297w485w490w496w(0) <= wire_addr_reg_w_lg_w_lg_w_q_range297w485w490w(0) AND wire_addr_reg_w_q_range495w(0);
	wire_addr_reg_w_lg_w_lg_w_q_range297w480w481w(0) <= wire_addr_reg_w_lg_w_q_range297w480w(0) AND bp1_wire;
	wire_addr_reg_w_lg_w_lg_w_q_range297w485w486w(0) <= wire_addr_reg_w_lg_w_q_range297w485w(0) AND bp2_wire;
	wire_addr_reg_w_lg_w_lg_w_q_range297w485w490w(0) <= wire_addr_reg_w_lg_w_q_range297w485w(0) AND wire_addr_reg_w_q_range489w(0);
	wire_addr_reg_w_lg_w_q_range297w480w(0) <= wire_addr_reg_w_q_range297w(0) AND bp2_wire;
	wire_addr_reg_w_lg_w_q_range297w485w(0) <= wire_addr_reg_w_q_range297w(0) AND wire_addr_reg_w_q_range484w(0);
	wire_addr_reg_w_q_range505w(0) <= addr_reg(18);
	wire_addr_reg_w_q_range500w(0) <= addr_reg(19);
	wire_addr_reg_w_q_range495w(0) <= addr_reg(20);
	wire_addr_reg_w_q_range489w(0) <= addr_reg(21);
	wire_addr_reg_w_q_range272w <= addr_reg(22 DOWNTO 0);
	wire_addr_reg_w_q_range484w(0) <= addr_reg(22);
	wire_addr_reg_w_q_range297w(0) <= addr_reg(23);
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_asmi_opcode_reg_ena(0) = '1') THEN asmi_opcode_reg(0) <= wire_asmi_opcode_reg_d(0);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_asmi_opcode_reg_ena(1) = '1') THEN asmi_opcode_reg(1) <= wire_asmi_opcode_reg_d(1);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_asmi_opcode_reg_ena(2) = '1') THEN asmi_opcode_reg(2) <= wire_asmi_opcode_reg_d(2);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_asmi_opcode_reg_ena(3) = '1') THEN asmi_opcode_reg(3) <= wire_asmi_opcode_reg_d(3);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_asmi_opcode_reg_ena(4) = '1') THEN asmi_opcode_reg(4) <= wire_asmi_opcode_reg_d(4);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_asmi_opcode_reg_ena(5) = '1') THEN asmi_opcode_reg(5) <= wire_asmi_opcode_reg_d(5);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_asmi_opcode_reg_ena(6) = '1') THEN asmi_opcode_reg(6) <= wire_asmi_opcode_reg_d(6);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_asmi_opcode_reg_ena(7) = '1') THEN asmi_opcode_reg(7) <= wire_asmi_opcode_reg_d(7);
			END IF;
		END IF;
	END PROCESS;
	wire_asmi_opcode_reg_d <= ( wire_w_lg_w177w178w & wire_w209w);
	loop28 : FOR i IN 0 TO 7 GENERATE
		wire_asmi_opcode_reg_ena(i) <= wire_w_lg_load_opcode211w(0);
	END GENERATE loop28;
	wire_asmi_opcode_reg_w_q_range129w <= asmi_opcode_reg(6 DOWNTO 0);
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '0' AND clkin_wire'event) THEN buf_empty_reg <= wire_cmpr5_aeb;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '0' AND clkin_wire'event) THEN busy_det_reg <= wire_w_lg_busy_wire1w(0);
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '0' AND clkin_wire'event) THEN clr_addmsb_reg <= ((wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range82w87w293w294w(0) OR wire_w_lg_w_lg_w_lg_do_read245w246w292w(0)) OR wire_w_lg_w_lg_w_lg_do_sec_erase289w290w291w(0));
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '1' AND clkin_wire'event) THEN clr_endrbyte_reg <= ((((wire_w_lg_do_read301w(0) AND (NOT wire_gen_cntr_q(2))) AND wire_gen_cntr_q(1)) AND wire_gen_cntr_q(0)) OR clr_read_wire);
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '0' AND clkin_wire'event) THEN clr_rdid_reg <= end_operation;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '0' AND clkin_wire'event) THEN clr_rdid_reg2 <= clr_rdid_reg;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '0' AND clkin_wire'event) THEN clr_read_reg <= ((end_operation OR do_read_sid) OR do_sec_prot);
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '0' AND clkin_wire'event) THEN clr_read_reg2 <= clr_read_reg;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '0' AND clkin_wire'event) THEN clr_rstat_reg <= ((end_operation OR do_read_sid) OR do_read);
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '0' AND clkin_wire'event) THEN clr_rstat_reg2 <= clr_rstat_reg;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '0' AND clkin_wire'event) THEN clr_write_reg <= ((((((wire_w_lg_w555w556w(0) OR wire_w_lg_do_write55w(0)) OR wire_w_lg_w_lg_w_lg_w_lg_do_write378w552w553w554w(0)) OR do_read_sid) OR do_sec_prot) OR do_read) OR do_fast_read);
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '0' AND clkin_wire'event) THEN clr_write_reg2 <= clr_write_reg;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '0' AND clkin_wire'event) THEN cnt_bfend_reg <= cnt_bfend_wire_in;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '0' AND clkin_wire'event) THEN do_wrmemadd_reg <= (wire_wrstage_cntr_q(1) AND wire_wrstage_cntr_q(0));
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, end_operation)
	BEGIN
		IF (end_operation = '1') THEN dvalid_reg <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_dvalid_reg_ena = '1') THEN dvalid_reg <= (end_read_byte AND end_one_cyc_pos);
			END IF;
		END IF;
	END PROCESS;
	wire_dvalid_reg_ena <= wire_w_lg_do_read301w(0);
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '0' AND clkin_wire'event) THEN dvalid_reg2 <= dvalid_reg;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '0' AND clkin_wire'event) THEN end1_cyc_reg <= end1_cyc_reg_in_wire;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '1' AND clkin_wire'event) THEN end1_cyc_reg2 <= end_one_cycle;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '0' AND clkin_wire'event) THEN end_op_hdlyreg <= end_operation;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '1' AND clkin_wire'event) THEN end_op_reg <= ((((((((((wire_stage_cntr_w_lg_w_q_range82w87w(0) AND ((wire_w_lg_w_lg_w_lg_w_lg_do_read245w246w247w248w(0) OR (do_read AND end_read)) OR (do_fast_read AND end_fast_read))) OR (wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range82w85w240w241w(0) AND wire_w_lg_do_polling239w(0))) OR (((wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range82w85w234w235w(0) AND wire_addbyte_cntr_q(2)) AND wire_addbyte_cntr_q(1)) AND wire_addbyte_cntr_q(0))) OR (wire_w_lg_w_lg_start_poll231w232w(0) AND wire_w_lg_st_busy_wire95w(0))) OR wire_stage_cntr_w_lg_w_lg_w_lg_w_lg_w_q_range82w83w84w229w230w(0)) OR wire_w_lg_w_lg_w_lg_do_write57w58w59w(0)) OR wire_w_lg_w_lg_do_write48w226w(0)) OR wire_w_lg_do_write55w(0)) OR wire_stage_cntr_w225w(0)) OR wire_stage_cntr_w_lg_w220w221w(0));
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, clr_write_wire)
	BEGIN
		IF (clr_write_wire = '1') THEN end_pgwrop_reg <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_end_pgwrop_reg_ena = '1') THEN end_pgwrop_reg <= buf_empty;
			END IF;
		END IF;
	END PROCESS;
	wire_end_pgwrop_reg_ena <= ((cnt_bfend_reg AND do_write) AND shift_pgwr_data);
	PROCESS (clkin_wire, clr_endrbyte_reg)
	BEGIN
		IF (clr_endrbyte_reg = '1') THEN end_rbyte_reg <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_end_rbyte_reg_ena = '1') THEN end_rbyte_reg <= wire_w_lg_w_lg_w_lg_do_read301w345w346w(0);
			END IF;
		END IF;
	END PROCESS;
	wire_end_rbyte_reg_ena <= (wire_gen_cntr_w_lg_w_q_range92w93w(0) AND wire_gen_cntr_q(0));
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '1' AND clkin_wire'event) THEN end_read_reg <= (((wire_w_lg_rden_wire360w(0) AND wire_w_lg_do_read301w(0)) AND data_valid_wire) AND end_read_byte);
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '0' AND clkin_wire'event) THEN ill_erase_reg <= illegal_erase_b4out_wire;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '0' AND clkin_wire'event) THEN ill_write_reg <= illegal_write_b4out_wire;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '0' AND clkin_wire'event) THEN max_cnt_reg <= wire_cmpr4_aeb;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '1' AND clkin_wire'event) THEN maxcnt_shift_reg <= (wire_w_lg_w_lg_reach_max_cnt453w454w(0) AND wire_w_lg_do_write378w(0));
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '0' AND clkin_wire'event) THEN maxcnt_shift_reg2 <= maxcnt_shift_reg;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, end_ophdly)
	BEGIN
		IF (end_ophdly = '1') THEN ncs_reg <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_ncs_reg_ena = '1') THEN ncs_reg <= '1';
			END IF;
		END IF;
	END PROCESS;
	wire_ncs_reg_ena <= (wire_stage_cntr_w_lg_w_lg_w_q_range82w83w84w(0) AND end_one_cyc_pos);
	wire_ncs_reg_w_lg_q262w(0) <= NOT ncs_reg;
	PROCESS (clkin_wire, clr_write_wire)
	BEGIN
		IF (clr_write_wire = '1') THEN pgwrbuf_dataout(0) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_pgwrbuf_dataout_ena(0) = '1') THEN pgwrbuf_dataout(0) <= wire_pgwrbuf_dataout_d(0);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, clr_write_wire)
	BEGIN
		IF (clr_write_wire = '1') THEN pgwrbuf_dataout(1) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_pgwrbuf_dataout_ena(1) = '1') THEN pgwrbuf_dataout(1) <= wire_pgwrbuf_dataout_d(1);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, clr_write_wire)
	BEGIN
		IF (clr_write_wire = '1') THEN pgwrbuf_dataout(2) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_pgwrbuf_dataout_ena(2) = '1') THEN pgwrbuf_dataout(2) <= wire_pgwrbuf_dataout_d(2);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, clr_write_wire)
	BEGIN
		IF (clr_write_wire = '1') THEN pgwrbuf_dataout(3) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_pgwrbuf_dataout_ena(3) = '1') THEN pgwrbuf_dataout(3) <= wire_pgwrbuf_dataout_d(3);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, clr_write_wire)
	BEGIN
		IF (clr_write_wire = '1') THEN pgwrbuf_dataout(4) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_pgwrbuf_dataout_ena(4) = '1') THEN pgwrbuf_dataout(4) <= wire_pgwrbuf_dataout_d(4);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, clr_write_wire)
	BEGIN
		IF (clr_write_wire = '1') THEN pgwrbuf_dataout(5) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_pgwrbuf_dataout_ena(5) = '1') THEN pgwrbuf_dataout(5) <= wire_pgwrbuf_dataout_d(5);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, clr_write_wire)
	BEGIN
		IF (clr_write_wire = '1') THEN pgwrbuf_dataout(6) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_pgwrbuf_dataout_ena(6) = '1') THEN pgwrbuf_dataout(6) <= wire_pgwrbuf_dataout_d(6);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, clr_write_wire)
	BEGIN
		IF (clr_write_wire = '1') THEN pgwrbuf_dataout(7) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_pgwrbuf_dataout_ena(7) = '1') THEN pgwrbuf_dataout(7) <= wire_pgwrbuf_dataout_d(7);
			END IF;
		END IF;
	END PROCESS;
	wire_pgwrbuf_dataout_d <= ( wire_w_lg_w_lg_read_bufdly411w412w & wire_w_lg_read_bufdly416w);
	loop29 : FOR i IN 0 TO 7 GENERATE
		wire_pgwrbuf_dataout_ena(i) <= wire_w_lg_read_bufdly406w(0);
	END GENERATE loop29;
	wire_pgwrbuf_dataout_w_q_range407w <= pgwrbuf_dataout(6 DOWNTO 0);
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (rdid_load = '1') THEN rdid_out_reg <= ( read_dout_reg(7 DOWNTO 0));
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '1' AND clkin_wire'event) THEN read_bufdly_reg <= read_buf;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_data_reg_ena(0) = '1') THEN read_data_reg(0) <= wire_read_data_reg_d(0);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_data_reg_ena(1) = '1') THEN read_data_reg(1) <= wire_read_data_reg_d(1);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_data_reg_ena(2) = '1') THEN read_data_reg(2) <= wire_read_data_reg_d(2);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_data_reg_ena(3) = '1') THEN read_data_reg(3) <= wire_read_data_reg_d(3);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_data_reg_ena(4) = '1') THEN read_data_reg(4) <= wire_read_data_reg_d(4);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_data_reg_ena(5) = '1') THEN read_data_reg(5) <= wire_read_data_reg_d(5);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_data_reg_ena(6) = '1') THEN read_data_reg(6) <= wire_read_data_reg_d(6);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_data_reg_ena(7) = '1') THEN read_data_reg(7) <= wire_read_data_reg_d(7);
			END IF;
		END IF;
	END PROCESS;
	wire_read_data_reg_d <= ( read_data_reg_in_wire(7 DOWNTO 0));
	loop30 : FOR i IN 0 TO 7 GENERATE
		wire_read_data_reg_ena(i) <= wire_w348w(0);
	END GENERATE loop30;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_read_dout_reg_ena(0) = '1') THEN read_dout_reg(0) <= wire_read_dout_reg_d(0);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_read_dout_reg_ena(1) = '1') THEN read_dout_reg(1) <= wire_read_dout_reg_d(1);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_read_dout_reg_ena(2) = '1') THEN read_dout_reg(2) <= wire_read_dout_reg_d(2);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_read_dout_reg_ena(3) = '1') THEN read_dout_reg(3) <= wire_read_dout_reg_d(3);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_read_dout_reg_ena(4) = '1') THEN read_dout_reg(4) <= wire_read_dout_reg_d(4);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_read_dout_reg_ena(5) = '1') THEN read_dout_reg(5) <= wire_read_dout_reg_d(5);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_read_dout_reg_ena(6) = '1') THEN read_dout_reg(6) <= wire_read_dout_reg_d(6);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_read_dout_reg_ena(7) = '1') THEN read_dout_reg(7) <= wire_read_dout_reg_d(7);
			END IF;
		END IF;
	END PROCESS;
	wire_read_dout_reg_d <= ( read_dout_reg(6 DOWNTO 0) & wire_w_lg_data0out_wire317w);
	loop31 : FOR i IN 0 TO 7 GENERATE
		wire_read_dout_reg_ena(i) <= wire_w_lg_w_lg_stage4_wire314w315w(0);
	END GENERATE loop31;
	PROCESS (clkin_wire, clr_rdid_wire)
	BEGIN
		IF (clr_rdid_wire = '1') THEN read_rdid_reg <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (busy_wire = '0') THEN read_rdid_reg <= read_rdid;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, clr_read_wire)
	BEGIN
		IF (clr_read_wire = '1') THEN read_reg <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_read_reg_ena = '1') THEN read_reg <= read;
			END IF;
		END IF;
	END PROCESS;
	wire_read_reg_ena <= (wire_w_lg_busy_wire1w(0) AND rden_wire);
	PROCESS (clkin_wire, clr_rstat_wire)
	BEGIN
		IF (clr_rstat_wire = '1') THEN read_status_reg <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (busy_wire = '0') THEN read_status_reg <= read_status;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, clr_write_wire)
	BEGIN
		IF (clr_write_wire = '1') THEN sec_erase_reg <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_sec_erase_reg_ena = '1') THEN sec_erase_reg <= sector_erase;
			END IF;
		END IF;
	END PROCESS;
	wire_sec_erase_reg_ena <= (wire_w_lg_busy_wire1w(0) AND wren_wire);
	PROCESS (clkin_wire, end_ophdly)
	BEGIN
		IF (end_ophdly = '1') THEN shftpgwr_data_reg <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN shftpgwr_data_reg <= ((wire_stage_cntr_w_lg_w_q_range82w87w(0) AND wire_wrstage_cntr_q(1)) AND wire_wrstage_cntr_q(0));
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '1' AND clkin_wire'event) THEN shift_op_reg <= wire_stage_cntr_w_lg_w_lg_w_q_range82w83w84w(0);
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '0' AND clkin_wire'event) THEN stage2_reg <= wire_stage_cntr_w_lg_w_lg_w_q_range82w83w84w(0);
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '1' AND clkin_wire'event) THEN stage3_dly_reg <= wire_stage_cntr_w_lg_w_q_range82w85w(0);
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '0' AND clkin_wire'event) THEN stage3_reg <= wire_stage_cntr_w_lg_w_q_range82w85w(0);
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '0' AND clkin_wire'event) THEN stage4_reg <= wire_stage_cntr_w_lg_w_q_range82w87w(0);
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, clr_write_wire)
	BEGIN
		IF (clr_write_wire = '1') THEN start_wrpoll_reg <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_start_wrpoll_reg_ena = '1') THEN start_wrpoll_reg <= wire_stage_cntr_w_lg_w_q_range82w85w(0);
			END IF;
		END IF;
	END PROCESS;
	wire_start_wrpoll_reg_ena <= ((do_write_rstat AND do_polling) AND end_one_cycle);
	PROCESS (clkin_wire, clr_write_wire)
	BEGIN
		IF (clr_write_wire = '1') THEN start_wrpoll_reg2 <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN start_wrpoll_reg2 <= start_wrpoll_reg;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, clr_rstat_wire)
	BEGIN
		IF (clr_rstat_wire = '1') THEN statreg_int(0) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_statreg_int_ena(0) = '1') THEN statreg_int(0) <= wire_statreg_int_d(0);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, clr_rstat_wire)
	BEGIN
		IF (clr_rstat_wire = '1') THEN statreg_int(1) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_statreg_int_ena(1) = '1') THEN statreg_int(1) <= wire_statreg_int_d(1);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, clr_rstat_wire)
	BEGIN
		IF (clr_rstat_wire = '1') THEN statreg_int(2) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_statreg_int_ena(2) = '1') THEN statreg_int(2) <= wire_statreg_int_d(2);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, clr_rstat_wire)
	BEGIN
		IF (clr_rstat_wire = '1') THEN statreg_int(3) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_statreg_int_ena(3) = '1') THEN statreg_int(3) <= wire_statreg_int_d(3);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, clr_rstat_wire)
	BEGIN
		IF (clr_rstat_wire = '1') THEN statreg_int(4) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_statreg_int_ena(4) = '1') THEN statreg_int(4) <= wire_statreg_int_d(4);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, clr_rstat_wire)
	BEGIN
		IF (clr_rstat_wire = '1') THEN statreg_int(5) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_statreg_int_ena(5) = '1') THEN statreg_int(5) <= wire_statreg_int_d(5);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, clr_rstat_wire)
	BEGIN
		IF (clr_rstat_wire = '1') THEN statreg_int(6) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_statreg_int_ena(6) = '1') THEN statreg_int(6) <= wire_statreg_int_d(6);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, clr_rstat_wire)
	BEGIN
		IF (clr_rstat_wire = '1') THEN statreg_int(7) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_statreg_int_ena(7) = '1') THEN statreg_int(7) <= wire_statreg_int_d(7);
			END IF;
		END IF;
	END PROCESS;
	wire_statreg_int_d <= ( read_dout_reg(7 DOWNTO 0));
	loop32 : FOR i IN 0 TO 7 GENERATE
		wire_statreg_int_ena(i) <= wire_w_lg_w_lg_end_operation391w392w(0);
	END GENERATE loop32;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_statreg_out_ena(0) = '1') THEN statreg_out(0) <= wire_statreg_out_d(0);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_statreg_out_ena(1) = '1') THEN statreg_out(1) <= wire_statreg_out_d(1);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_statreg_out_ena(2) = '1') THEN statreg_out(2) <= wire_statreg_out_d(2);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_statreg_out_ena(3) = '1') THEN statreg_out(3) <= wire_statreg_out_d(3);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_statreg_out_ena(4) = '1') THEN statreg_out(4) <= wire_statreg_out_d(4);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_statreg_out_ena(5) = '1') THEN statreg_out(5) <= wire_statreg_out_d(5);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_statreg_out_ena(6) = '1') THEN statreg_out(6) <= wire_statreg_out_d(6);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire)
	BEGIN
		IF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_statreg_out_ena(7) = '1') THEN statreg_out(7) <= wire_statreg_out_d(7);
			END IF;
		END IF;
	END PROCESS;
	wire_statreg_out_d <= ( read_dout_reg(7 DOWNTO 0));
	loop33 : FOR i IN 0 TO 7 GENERATE
		wire_statreg_out_ena(i) <= wire_w383w(0);
	END GENERATE loop33;
	PROCESS (clkin_wire, clr_write_wire)
	BEGIN
		IF (clr_write_wire = '1') THEN write_prot_reg <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_write_prot_reg_ena = '1') THEN write_prot_reg <= ((wire_w_lg_do_write57w(0) AND ((((((wire_addr_reg_w_lg_w_lg_w_lg_w506w507w508w509w(0) OR (wire_addr_reg_w_lg_w502w503w(0) AND wire_w_lg_bp0_wire479w(0))) OR wire_addr_reg_w_lg_w498w499w(0)) OR ((wire_addr_reg_w_lg_w_lg_w_lg_w_q_range297w485w490w491w(0) AND wire_w_lg_bp1_wire483w(0)) AND wire_w_lg_bp0_wire479w(0))) OR wire_addr_reg_w_lg_w_lg_w_lg_w_lg_w_q_range297w485w486w487w488w(0)) OR (wire_addr_reg_w_lg_w_lg_w_q_range297w480w481w(0) AND wire_w_lg_bp0_wire479w(0))) OR wire_w_lg_w_lg_bp2_wire477w478w(0))) OR be_write_prot);
			END IF;
		END IF;
	END PROCESS;
	wire_write_prot_reg_ena <= (((wire_w_lg_w_lg_do_sec_erase468w469w(0) AND (NOT wire_wrstage_cntr_q(1))) AND wire_wrstage_cntr_q(0)) AND end_ophdly);
	PROCESS (clkin_wire, clr_write_wire)
	BEGIN
		IF (clr_write_wire = '1') THEN write_reg <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_write_reg_ena = '1') THEN write_reg <= write;
			END IF;
		END IF;
	END PROCESS;
	wire_write_reg_ena <= (wire_w_lg_busy_wire1w(0) AND wren_wire);
	PROCESS (clkin_wire, clr_write_wire)
	BEGIN
		IF (clr_write_wire = '1') THEN write_rstat_reg <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN write_rstat_reg <= (wire_w_lg_w_lg_do_write57w58w(0) AND (((NOT wire_wrstage_cntr_q(1)) AND wire_wrstage_cntr_w_lg_w_q_range460w461w(0)) OR wire_wrstage_cntr_w_lg_w_q_range462w463w(0)));
		END IF;
	END PROCESS;
	wire_cmpr4_dataa <= ( page_size_wire(8 DOWNTO 0));
	wire_cmpr4_datab <= ( wire_pgwr_data_cntr_q(8 DOWNTO 0));
	cmpr4 :  lpm_compare
	  GENERIC MAP (
		LPM_WIDTH => 9
	  )
	  PORT MAP ( 
		aeb => wire_cmpr4_aeb,
		dataa => wire_cmpr4_dataa,
		datab => wire_cmpr4_datab
	  );
	wire_cmpr5_dataa <= ( wire_pgwr_data_cntr_q(8 DOWNTO 0));
	wire_cmpr5_datab <= ( wire_pgwr_read_cntr_q(8 DOWNTO 0));
	cmpr5 :  lpm_compare
	  GENERIC MAP (
		LPM_WIDTH => 9
	  )
	  PORT MAP ( 
		aeb => wire_cmpr5_aeb,
		dataa => wire_cmpr5_dataa,
		datab => wire_cmpr5_datab
	  );
	wire_pgwr_data_cntr_clk_en <= wire_w_lg_w_lg_w_lg_shift_bytes_wire403w419w420w(0);
	wire_w_lg_w_lg_w_lg_shift_bytes_wire403w419w420w(0) <= ((shift_bytes_wire AND wren_wire) AND wire_w_lg_reach_max_cnt418w(0)) AND wire_w_lg_do_write378w(0);
	wire_pgwr_data_cntr_w_q_range424w(0) <= wire_pgwr_data_cntr_q(1);
	wire_pgwr_data_cntr_w_q_range427w(0) <= wire_pgwr_data_cntr_q(2);
	wire_pgwr_data_cntr_w_q_range430w(0) <= wire_pgwr_data_cntr_q(3);
	wire_pgwr_data_cntr_w_q_range433w(0) <= wire_pgwr_data_cntr_q(4);
	wire_pgwr_data_cntr_w_q_range436w(0) <= wire_pgwr_data_cntr_q(5);
	wire_pgwr_data_cntr_w_q_range439w(0) <= wire_pgwr_data_cntr_q(6);
	wire_pgwr_data_cntr_w_q_range442w(0) <= wire_pgwr_data_cntr_q(7);
	wire_pgwr_data_cntr_w_q_range445w(0) <= wire_pgwr_data_cntr_q(8);
	pgwr_data_cntr :  lpm_counter
	  GENERIC MAP (
		lpm_direction => "UP",
		lpm_port_updown => "PORT_UNUSED",
		lpm_width => 9
	  )
	  PORT MAP ( 
		aclr => clr_write_wire,
		clk_en => wire_pgwr_data_cntr_clk_en,
		clock => clkin_wire,
		q => wire_pgwr_data_cntr_q
	  );
	pgwr_read_cntr :  lpm_counter
	  GENERIC MAP (
		lpm_direction => "UP",
		lpm_port_updown => "PORT_UNUSED",
		lpm_width => 9
	  )
	  PORT MAP ( 
		aclr => clr_write_wire,
		clk_en => read_buf,
		clock => clkin_wire,
		q => wire_pgwr_read_cntr_q
	  );
	wire_mux211_dataout <= end_add_cycle_mux_datab_wire WHEN do_fast_read = '1'  ELSE wire_addbyte_cntr_w_lg_w_q_range123w124w(0);
	wire_scfifo3_data <= ( datain(7 DOWNTO 0));
	wire_scfifo3_rdreq <= wire_w_lg_read_buf405w(0);
	wire_w_lg_read_buf405w(0) <= read_buf OR dummy_read_buf;
	wire_scfifo3_wrreq <= wire_w_lg_w_lg_shift_bytes_wire403w404w(0);
	wire_w_lg_w_lg_shift_bytes_wire403w404w(0) <= (shift_bytes_wire AND wren_wire) AND wire_w_lg_do_write378w(0);
	wire_scfifo3_w_q_range410w <= wire_scfifo3_q(7 DOWNTO 1);
	wire_scfifo3_w_q_range415w(0) <= wire_scfifo3_q(0);
	scfifo3 :  scfifo
	  GENERIC MAP (
		LPM_NUMWORDS => 258,
		LPM_WIDTH => 8,
		LPM_WIDTHU => 9,
		USE_EAB => "ON"
	  )
	  PORT MAP ( 
		aclr => clr_write_wire,
		clock => clkin_wire,
		data => wire_scfifo3_data,
		q => wire_scfifo3_q,
		rdreq => wire_scfifo3_rdreq,
		wrreq => wire_scfifo3_wrreq
	  );
	stratixii_asmiblock2 :  arriaii_asmiblock
	  PORT MAP ( 
		data0out => wire_stratixii_asmiblock2_data0out,
		dclkin => clkin_wire,
		oe => oe_wire,
		scein => scein_wire,
		sdoin => sdoin_wire
	  );

 END RTL; --flash_access_altasmi_parallel_era2
--VALID FILE


LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY flash_access IS
	PORT
	(
		addr		: IN STD_LOGIC_VECTOR (23 DOWNTO 0);
		clkin		: IN STD_LOGIC ;
		datain		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		rden		: IN STD_LOGIC ;
		read		: IN STD_LOGIC ;
		read_rdid		: IN STD_LOGIC ;
		read_status		: IN STD_LOGIC ;
		sector_erase		: IN STD_LOGIC ;
		shift_bytes		: IN STD_LOGIC ;
		wren		: IN STD_LOGIC ;
		write		: IN STD_LOGIC ;
		busy		: OUT STD_LOGIC ;
		data_valid		: OUT STD_LOGIC ;
		dataout		: OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
		illegal_erase		: OUT STD_LOGIC ;
		illegal_write		: OUT STD_LOGIC ;
		rdid_out		: OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
		status_out		: OUT STD_LOGIC_VECTOR (7 DOWNTO 0)
	);
END flash_access;


ARCHITECTURE RTL OF flash_access IS

	ATTRIBUTE synthesis_clearbox: natural;
	ATTRIBUTE synthesis_clearbox OF RTL: ARCHITECTURE IS 2;
	ATTRIBUTE clearbox_macroname: string;
	ATTRIBUTE clearbox_macroname OF RTL: ARCHITECTURE IS "ALTASMI_PARALLEL";
	ATTRIBUTE clearbox_defparam: string;
	ATTRIBUTE clearbox_defparam OF RTL: ARCHITECTURE IS "data_width=STANDARD;epcs_type=EPCS128;intended_device_family=Arria II GX;lpm_hint=UNUSED;lpm_type=altasmi_parallel;page_size=256;port_bulk_erase=PORT_UNUSED;port_fast_read=PORT_UNUSED;port_illegal_erase=PORT_USED;port_illegal_write=PORT_USED;port_rdid_out=PORT_USED;port_read_address=PORT_UNUSED;port_read_rdid=PORT_USED;port_read_sid=PORT_UNUSED;port_read_status=PORT_USED;port_sector_erase=PORT_USED;port_sector_protect=PORT_UNUSED;port_shift_bytes=PORT_USED;port_wren=PORT_USED;port_write=PORT_USED;use_eab=ON;";
	SIGNAL sub_wire0	: STD_LOGIC ;
	SIGNAL sub_wire1	: STD_LOGIC ;
	SIGNAL sub_wire2	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire3	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire4	: STD_LOGIC ;
	SIGNAL sub_wire5	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire6	: STD_LOGIC ;



	COMPONENT flash_access_altasmi_parallel_era2
	PORT (
			clkin	: IN STD_LOGIC ;
			data_valid	: OUT STD_LOGIC ;
			datain	: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
			illegal_erase	: OUT STD_LOGIC ;
			rden	: IN STD_LOGIC ;
			dataout	: OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
			rdid_out	: OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
			read_rdid	: IN STD_LOGIC ;
			addr	: IN STD_LOGIC_VECTOR (23 DOWNTO 0);
			busy	: OUT STD_LOGIC ;
			read_status	: IN STD_LOGIC ;
			sector_erase	: IN STD_LOGIC ;
			status_out	: OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
			write	: IN STD_LOGIC ;
			illegal_write	: OUT STD_LOGIC ;
			read	: IN STD_LOGIC ;
			shift_bytes	: IN STD_LOGIC ;
			wren	: IN STD_LOGIC 
	);
	END COMPONENT;

BEGIN
	data_valid    <= sub_wire0;
	illegal_erase    <= sub_wire1;
	dataout    <= sub_wire2(7 DOWNTO 0);
	rdid_out    <= sub_wire3(7 DOWNTO 0);
	busy    <= sub_wire4;
	status_out    <= sub_wire5(7 DOWNTO 0);
	illegal_write    <= sub_wire6;

	flash_access_altasmi_parallel_era2_component : flash_access_altasmi_parallel_era2
	PORT MAP (
		clkin => clkin,
		datain => datain,
		rden => rden,
		read_rdid => read_rdid,
		addr => addr,
		read_status => read_status,
		sector_erase => sector_erase,
		write => write,
		read => read,
		shift_bytes => shift_bytes,
		wren => wren,
		data_valid => sub_wire0,
		illegal_erase => sub_wire1,
		dataout => sub_wire2,
		rdid_out => sub_wire3,
		busy => sub_wire4,
		status_out => sub_wire5,
		illegal_write => sub_wire6
	);



END RTL;

-- ============================================================
-- CNX file retrieval info
-- ============================================================
-- Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
-- Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Arria II GX"
-- Retrieval info: CONSTANT: DATA_WIDTH STRING "STANDARD"
-- Retrieval info: CONSTANT: EPCS_TYPE STRING "EPCS128"
-- Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "Arria II GX"
-- Retrieval info: CONSTANT: LPM_HINT STRING "UNUSED"
-- Retrieval info: CONSTANT: LPM_TYPE STRING "altasmi_parallel"
-- Retrieval info: CONSTANT: PAGE_SIZE NUMERIC "256"
-- Retrieval info: CONSTANT: PORT_BULK_ERASE STRING "PORT_UNUSED"
-- Retrieval info: CONSTANT: PORT_FAST_READ STRING "PORT_UNUSED"
-- Retrieval info: CONSTANT: PORT_ILLEGAL_ERASE STRING "PORT_USED"
-- Retrieval info: CONSTANT: PORT_ILLEGAL_WRITE STRING "PORT_USED"
-- Retrieval info: CONSTANT: PORT_RDID_OUT STRING "PORT_USED"
-- Retrieval info: CONSTANT: PORT_READ_ADDRESS STRING "PORT_UNUSED"
-- Retrieval info: CONSTANT: PORT_READ_RDID STRING "PORT_USED"
-- Retrieval info: CONSTANT: PORT_READ_SID STRING "PORT_UNUSED"
-- Retrieval info: CONSTANT: PORT_READ_STATUS STRING "PORT_USED"
-- Retrieval info: CONSTANT: PORT_SECTOR_ERASE STRING "PORT_USED"
-- Retrieval info: CONSTANT: PORT_SECTOR_PROTECT STRING "PORT_UNUSED"
-- Retrieval info: CONSTANT: PORT_SHIFT_BYTES STRING "PORT_USED"
-- Retrieval info: CONSTANT: PORT_WREN STRING "PORT_USED"
-- Retrieval info: CONSTANT: PORT_WRITE STRING "PORT_USED"
-- Retrieval info: CONSTANT: USE_EAB STRING "ON"
-- Retrieval info: USED_PORT: addr 0 0 24 0 INPUT NODEFVAL "addr[23..0]"
-- Retrieval info: CONNECT: @addr 0 0 24 0 addr 0 0 24 0
-- Retrieval info: USED_PORT: busy 0 0 0 0 OUTPUT NODEFVAL "busy"
-- Retrieval info: CONNECT: busy 0 0 0 0 @busy 0 0 0 0
-- Retrieval info: USED_PORT: clkin 0 0 0 0 INPUT NODEFVAL "clkin"
-- Retrieval info: CONNECT: @clkin 0 0 0 0 clkin 0 0 0 0
-- Retrieval info: USED_PORT: data_valid 0 0 0 0 OUTPUT NODEFVAL "data_valid"
-- Retrieval info: CONNECT: data_valid 0 0 0 0 @data_valid 0 0 0 0
-- Retrieval info: USED_PORT: datain 0 0 8 0 INPUT NODEFVAL "datain[7..0]"
-- Retrieval info: CONNECT: @datain 0 0 8 0 datain 0 0 8 0
-- Retrieval info: USED_PORT: dataout 0 0 8 0 OUTPUT NODEFVAL "dataout[7..0]"
-- Retrieval info: CONNECT: dataout 0 0 8 0 @dataout 0 0 8 0
-- Retrieval info: USED_PORT: illegal_erase 0 0 0 0 OUTPUT NODEFVAL "illegal_erase"
-- Retrieval info: CONNECT: illegal_erase 0 0 0 0 @illegal_erase 0 0 0 0
-- Retrieval info: USED_PORT: illegal_write 0 0 0 0 OUTPUT NODEFVAL "illegal_write"
-- Retrieval info: CONNECT: illegal_write 0 0 0 0 @illegal_write 0 0 0 0
-- Retrieval info: USED_PORT: rden 0 0 0 0 INPUT NODEFVAL "rden"
-- Retrieval info: CONNECT: @rden 0 0 0 0 rden 0 0 0 0
-- Retrieval info: USED_PORT: rdid_out 0 0 8 0 OUTPUT NODEFVAL "rdid_out[7..0]"
-- Retrieval info: CONNECT: rdid_out 0 0 8 0 @rdid_out 0 0 8 0
-- Retrieval info: USED_PORT: read 0 0 0 0 INPUT NODEFVAL "read"
-- Retrieval info: CONNECT: @read 0 0 0 0 read 0 0 0 0
-- Retrieval info: USED_PORT: read_rdid 0 0 0 0 INPUT NODEFVAL "read_rdid"
-- Retrieval info: CONNECT: @read_rdid 0 0 0 0 read_rdid 0 0 0 0
-- Retrieval info: USED_PORT: read_status 0 0 0 0 INPUT NODEFVAL "read_status"
-- Retrieval info: CONNECT: @read_status 0 0 0 0 read_status 0 0 0 0
-- Retrieval info: USED_PORT: sector_erase 0 0 0 0 INPUT NODEFVAL "sector_erase"
-- Retrieval info: CONNECT: @sector_erase 0 0 0 0 sector_erase 0 0 0 0
-- Retrieval info: USED_PORT: shift_bytes 0 0 0 0 INPUT NODEFVAL "shift_bytes"
-- Retrieval info: CONNECT: @shift_bytes 0 0 0 0 shift_bytes 0 0 0 0
-- Retrieval info: USED_PORT: status_out 0 0 8 0 OUTPUT NODEFVAL "status_out[7..0]"
-- Retrieval info: CONNECT: status_out 0 0 8 0 @status_out 0 0 8 0
-- Retrieval info: USED_PORT: wren 0 0 0 0 INPUT NODEFVAL "wren"
-- Retrieval info: CONNECT: @wren 0 0 0 0 wren 0 0 0 0
-- Retrieval info: USED_PORT: write 0 0 0 0 INPUT NODEFVAL "write"
-- Retrieval info: CONNECT: @write 0 0 0 0 write 0 0 0 0
-- Retrieval info: GEN_FILE: TYPE_NORMAL flash_access.vhd TRUE FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL flash_access.qip TRUE FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL flash_access.bsf TRUE TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL flash_access_inst.vhd TRUE TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL flash_access.inc TRUE TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL flash_access.cmp TRUE TRUE
